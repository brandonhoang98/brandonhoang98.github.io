// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/VCC.v,v 1.8 2003/01/21 01:55:44 wloo Exp $

/*

FUNCTION	: VCC cell

*/

`timescale  100 ps / 10 ps


module VCC(P);

    output P;

	assign P = 1'b1;

endmodule

