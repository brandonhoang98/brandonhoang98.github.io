// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/PPC405.v,v 1.10 2003/01/21 01:55:40 wloo Exp $

/*

		: Power PC

*/

`timescale  1 ps / 1 ps

module PPC405 (
		C405CPMCORESLEEPREQ,
		C405CPMMSRCE,
		C405CPMMSREE,
		C405CPMTIMERIRQ,
		C405CPMTIMERRESETREQ,
		C405DBGMSRWE,
		C405DBGSTOPACK,
		C405DBGWBCOMPLETE,
		C405DBGWBFULL,
		C405DBGWBIAR,
		C405DCRABUS,
		C405DCRDBUSOUT,
		C405DCRREAD,
		C405DCRWRITE,
		C405JTGCAPTUREDR,
		C405JTGEXTEST,
		C405JTGPGMOUT,
		C405JTGSHIFTDR,
		C405JTGTDO,
		C405JTGTDOEN,
		C405JTGUPDATEDR,
		C405PLBDCUABORT,
		C405PLBDCUABUS,
		C405PLBDCUBE,
		C405PLBDCUCACHEABLE,
		C405PLBDCUGUARDED,
		C405PLBDCUPRIORITY,
		C405PLBDCUREQUEST,
		C405PLBDCURNW,
		C405PLBDCUSIZE2,
		C405PLBDCUU0ATTR,
		C405PLBDCUWRDBUS,
		C405PLBDCUWRITETHRU,
		C405PLBICUABORT,
		C405PLBICUABUS,
		C405PLBICUCACHEABLE,
		C405PLBICUPRIORITY,
		C405PLBICUREQUEST,
		C405PLBICUSIZE,
		C405PLBICUU0ATTR,
		C405RSTCHIPRESETREQ,
		C405RSTCORERESETREQ,
		C405RSTSYSRESETREQ,
		C405TRCCYCLE,
		C405TRCEVENEXECUTIONSTATUS,
		C405TRCODDEXECUTIONSTATUS,
		C405TRCTRACESTATUS,
		C405TRCTRIGGEREVENTOUT,
		C405TRCTRIGGEREVENTTYPE,
		C405XXXMACHINECHECK,
		DSOCMBRAMABUS,
		DSOCMBRAMBYTEWRITE,
		DSOCMBRAMEN,
		DSOCMBRAMWRDBUS,
		DSOCMBUSY,
		ISOCMBRAMEN,
		ISOCMBRAMEVENWRITEEN,
		ISOCMBRAMODDWRITEEN,
		ISOCMBRAMRDABUS,
		ISOCMBRAMWRABUS,
		ISOCMBRAMWRDBUS,

		BRAMDSOCMCLK,
		BRAMDSOCMRDDBUS,
		BRAMISOCMCLK,
		BRAMISOCMRDDBUS,
		CPMC405CLOCK,
		CPMC405CORECLKINACTIVE,
		CPMC405CPUCLKEN,
		CPMC405JTAGCLKEN,
		CPMC405TIMERCLKEN,
		CPMC405TIMERTICK,
		DBGC405DEBUGHALT,
		DBGC405EXTBUSHOLDACK,
		DBGC405UNCONDDEBUGEVENT,
		DCRC405ACK,
		DCRC405DBUSIN,
		DSARCVALUE,
		DSCNTLVALUE,
		EICC405CRITINPUTIRQ,
		EICC405EXTINPUTIRQ,
		ISARCVALUE,
		ISCNTLVALUE,
		JTGC405BNDSCANTDO,
		JTGC405TCK,
		JTGC405TDI,
		JTGC405TMS,
		JTGC405TRSTNEG,
		MCBCPUCLKEN,
		MCBJTAGEN,
		MCBTIMEREN,
		MCPPCRST,
		PLBC405DCUADDRACK,
		PLBC405DCUBUSY,
		PLBC405DCUERR,
		PLBC405DCURDDACK,
		PLBC405DCURDDBUS,
		PLBC405DCURDWDADDR,
		PLBC405DCUSSIZE1,
		PLBC405DCUWRDACK,
		PLBC405ICUADDRACK,
		PLBC405ICUBUSY,
		PLBC405ICUERR,
		PLBC405ICURDDACK,
		PLBC405ICURDDBUS,
		PLBC405ICURDWDADDR,
		PLBC405ICUSSIZE1,
		PLBCLK,
		RSTC405RESETCHIP,
		RSTC405RESETCORE,
		RSTC405RESETSYS,
		TIEC405DETERMINISTICMULT,
		TIEC405DISOPERANDFWD,
		TIEC405MMUEN,
		TIEDSOCMDCRADDR,
		TIEISOCMDCRADDR,
		TRCC405TRACEDISABLE,
		TRCC405TRIGGEREVENTIN
);

parameter in_delay=10;
parameter out_delay=10;
parameter PPCUSER = 4'b0000;

output		C405CPMCORESLEEPREQ;
output		C405CPMMSRCE;
output		C405CPMMSREE;
output		C405CPMTIMERIRQ;
output		C405CPMTIMERRESETREQ;
output		C405DBGMSRWE;
output		C405DBGSTOPACK;
output		C405DBGWBCOMPLETE;
output		C405DBGWBFULL;
output	[0:29]	C405DBGWBIAR;
output	[0:9]	C405DCRABUS;
output	[0:31]	C405DCRDBUSOUT;
output		C405DCRREAD;
output		C405DCRWRITE;
output		C405JTGCAPTUREDR;
output		C405JTGEXTEST;
output		C405JTGPGMOUT;
output		C405JTGSHIFTDR;
output		C405JTGTDO;
output		C405JTGTDOEN;
output		C405JTGUPDATEDR;
output		C405PLBDCUABORT;
output	[0:31]	C405PLBDCUABUS;
output	[0:7]	C405PLBDCUBE;
output		C405PLBDCUCACHEABLE;
output		C405PLBDCUGUARDED;
output	[0:1]	C405PLBDCUPRIORITY;
output		C405PLBDCUREQUEST;
output		C405PLBDCURNW;
output		C405PLBDCUSIZE2;
output		C405PLBDCUU0ATTR;
output	[0:63]	C405PLBDCUWRDBUS;
output		C405PLBDCUWRITETHRU;
output		C405PLBICUABORT;
output	[0:29]	C405PLBICUABUS;
output		C405PLBICUCACHEABLE;
output	[0:1]	C405PLBICUPRIORITY;
output		C405PLBICUREQUEST;
output	[2:3]	C405PLBICUSIZE;
output		C405PLBICUU0ATTR;
output		C405RSTCHIPRESETREQ;
output		C405RSTCORERESETREQ;
output		C405RSTSYSRESETREQ;
output		C405TRCCYCLE;
output	[0:1]	C405TRCEVENEXECUTIONSTATUS;
output	[0:1]	C405TRCODDEXECUTIONSTATUS;
output	[0:3]	C405TRCTRACESTATUS;
output		C405TRCTRIGGEREVENTOUT;
output	[0:10]	C405TRCTRIGGEREVENTTYPE;
output		C405XXXMACHINECHECK;
output	[8:29]	DSOCMBRAMABUS;
output	[0:3]	DSOCMBRAMBYTEWRITE;
output		DSOCMBRAMEN;
output	[0:31]	DSOCMBRAMWRDBUS;
output		DSOCMBUSY;
output		ISOCMBRAMEN;
output		ISOCMBRAMEVENWRITEEN;
output		ISOCMBRAMODDWRITEEN;
output	[8:28]	ISOCMBRAMRDABUS;
output	[8:28]	ISOCMBRAMWRABUS;
output	[0:31]	ISOCMBRAMWRDBUS;

input		BRAMDSOCMCLK;
input	[0:31]	BRAMDSOCMRDDBUS;
input		BRAMISOCMCLK;
input	[0:63]	BRAMISOCMRDDBUS;
input		CPMC405CLOCK;
input		CPMC405CORECLKINACTIVE;
input		CPMC405CPUCLKEN;
input		CPMC405JTAGCLKEN;
input		CPMC405TIMERCLKEN;
input		CPMC405TIMERTICK;
input		DBGC405DEBUGHALT;
input		DBGC405EXTBUSHOLDACK;
input		DBGC405UNCONDDEBUGEVENT;
input		DCRC405ACK;
input	[0:31]	DCRC405DBUSIN;
input	[0:7]	DSARCVALUE;
input	[0:7]	DSCNTLVALUE;
input		EICC405CRITINPUTIRQ;
input		EICC405EXTINPUTIRQ;
input	[0:7]	ISARCVALUE;
input	[0:7]	ISCNTLVALUE;
input		JTGC405BNDSCANTDO;
input		JTGC405TCK;
input		JTGC405TDI;
input		JTGC405TMS;
input		JTGC405TRSTNEG;
input		MCBCPUCLKEN;
input		MCBJTAGEN;
input		MCBTIMEREN;
input		MCPPCRST;
input		PLBC405DCUADDRACK;
input		PLBC405DCUBUSY;
input		PLBC405DCUERR;
input		PLBC405DCURDDACK;
input	[0:63]	PLBC405DCURDDBUS;
input	[1:3]	PLBC405DCURDWDADDR;
input		PLBC405DCUSSIZE1;
input		PLBC405DCUWRDACK;
input		PLBC405ICUADDRACK;
input		PLBC405ICUBUSY;
input		PLBC405ICUERR;
input		PLBC405ICURDDACK;
input	[0:63]	PLBC405ICURDDBUS;
input	[1:3]	PLBC405ICURDWDADDR;
input		PLBC405ICUSSIZE1;
input		PLBCLK;
input		RSTC405RESETCHIP;
input		RSTC405RESETCORE;
input		RSTC405RESETSYS;
input		TIEC405DETERMINISTICMULT;
input		TIEC405DISOPERANDFWD;
input		TIEC405MMUEN;
input	[0:7]	TIEDSOCMDCRADDR;
input	[0:7]	TIEISOCMDCRADDR;
input		TRCC405TRACEDISABLE;
input		TRCC405TRIGGEREVENTIN;

// define input delay bus

wire [0:31] BRAMDSOCMRDDBUS_delay;
wire [0:63] BRAMISOCMRDDBUS_delay;
wire [0:31] DCRC405DBUSIN_delay;
wire [0:7] DSARCVALUE_delay;
wire [0:7] DSCNTLVALUE_delay;
wire [0:7] ISARCVALUE_delay;
wire [0:7] ISCNTLVALUE_delay;
wire [0:63] PLBC405DCURDDBUS_delay;
wire [1:3] PLBC405DCURDWDADDR_delay;
wire [0:63] PLBC405ICURDDBUS_delay;
wire [1:3] PLBC405ICURDWDADDR_delay;
wire [0:7] TIEDSOCMDCRADDR_delay;
wire [0:7] TIEISOCMDCRADDR_delay;

// define input delay pins

wire CPMC405CORECLKINACTIVE_delay;
wire CPMC405CPUCLKEN_delay;
wire CPMC405JTAGCLKEN_delay;
wire CPMC405TIMERCLKEN_delay;
wire CPMC405TIMERTICK_delay;
wire DBGC405DEBUGHALT_delay;
wire DBGC405EXTBUSHOLDACK_delay;
wire DBGC405UNCONDDEBUGEVENT_delay;
wire DCRC405ACK_delay;
wire EICC405CRITINPUTIRQ_delay;
wire EICC405EXTINPUTIRQ_delay;
wire JTGC405BNDSCANTDO_delay;
wire JTGC405TCK_delay;
wire JTGC405TDI_delay;
wire JTGC405TMS_delay;
wire JTGC405TRSTNEG_delay;
wire MCBCPUCLKEN_delay;
wire MCBJTAGEN_delay;
wire MCBTIMEREN_delay;
wire MCPPCRST_delay;
wire PLBC405DCUADDRACK_delay;
wire PLBC405DCUBUSY_delay;
wire PLBC405DCUERR_delay;
wire PLBC405DCURDDACK_delay;
wire PLBC405DCUSSIZE1_delay;
wire PLBC405DCUWRDACK_delay;
wire PLBC405ICUADDRACK_delay;
wire PLBC405ICUBUSY_delay;
wire PLBC405ICUERR_delay;
wire PLBC405ICURDDACK_delay;
wire PLBC405ICUSSIZE1_delay;
wire RSTC405RESETCHIP_delay;
wire RSTC405RESETCORE_delay;
wire RSTC405RESETSYS_delay;
wire TIEC405DETERMINISTICMULT_delay;
wire TIEC405DISOPERANDFWD_delay;
wire TIEC405MMUEN_delay;
wire TRCC405TRACEDISABLE_delay;
wire TRCC405TRIGGEREVENTIN_delay;

// define output delay bus

wire [0:29] C405DBGWBIAR_delay;
wire [0:9] C405DCRABUS_delay;
wire [0:31] C405DCRDBUSOUT_delay;
wire [0:31] C405PLBDCUABUS_delay;
wire [0:7] C405PLBDCUBE_delay;
wire [0:1] C405PLBDCUPRIORITY_delay;
wire [0:63] C405PLBDCUWRDBUS_delay;
wire [0:29] C405PLBICUABUS_delay;
wire [0:1] C405PLBICUPRIORITY_delay;
wire [2:3] C405PLBICUSIZE_delay;
wire [0:1] C405TRCEVENEXECUTIONSTATUS_delay;
wire [0:1] C405TRCODDEXECUTIONSTATUS_delay;
wire [0:3] C405TRCTRACESTATUS_delay;
wire [0:10] C405TRCTRIGGEREVENTTYPE_delay;
wire [8:29] DSOCMBRAMABUS_delay;
wire [0:3] DSOCMBRAMBYTEWRITE_delay;
wire [0:31] DSOCMBRAMWRDBUS_delay;
wire [8:28] ISOCMBRAMRDABUS_delay;
wire [8:28] ISOCMBRAMWRABUS_delay;
wire [0:31] ISOCMBRAMWRDBUS_delay;

// define output delay pins

wire C405CPMCORESLEEPREQ_delay;
wire C405CPMMSRCE_delay;
wire C405CPMMSREE_delay;
wire C405CPMTIMERIRQ_delay;
wire C405CPMTIMERRESETREQ_delay;
wire C405DBGMSRWE_delay;
wire C405DBGSTOPACK_delay;
wire C405DBGWBCOMPLETE_delay;
wire C405DBGWBFULL_delay;
wire C405DCRREAD_delay;
wire C405DCRWRITE_delay;
wire C405JTGCAPTUREDR_delay;
wire C405JTGEXTEST_delay;
wire C405JTGPGMOUT_delay;
wire C405JTGSHIFTDR_delay;
wire C405JTGTDO_delay;
wire C405JTGTDOEN_delay;
wire C405JTGUPDATEDR_delay;
wire C405PLBDCUABORT_delay;
wire C405PLBDCUCACHEABLE_delay;
wire C405PLBDCUGUARDED_delay;
wire C405PLBDCUREQUEST_delay;
wire C405PLBDCURNW_delay;
wire C405PLBDCUSIZE2_delay;
wire C405PLBDCUU0ATTR_delay;
wire C405PLBDCUWRITETHRU_delay;
wire C405PLBICUABORT_delay;
wire C405PLBICUCACHEABLE_delay;
wire C405PLBICUREQUEST_delay;
wire C405PLBICUU0ATTR_delay;
wire C405RSTCHIPRESETREQ_delay;
wire C405RSTCORERESETREQ_delay;
wire C405RSTSYSRESETREQ_delay;
wire C405TRCCYCLE_delay;
wire C405TRCTRIGGEREVENTOUT_delay;
wire C405XXXMACHINECHECK_delay;
wire DSOCMBRAMEN_delay;
wire DSOCMBUSY_delay;
wire ISOCMBRAMEN_delay;
wire ISOCMBRAMEVENWRITEEN_delay;
wire ISOCMBRAMODDWRITEEN_delay;

assign #(in_delay) BRAMDSOCMRDDBUS_delay[0:31] = BRAMDSOCMRDDBUS[0:31];
assign #(in_delay) BRAMISOCMRDDBUS_delay[0:63] = BRAMISOCMRDDBUS[0:63];
assign #(in_delay) CPMC405CORECLKINACTIVE_delay = CPMC405CORECLKINACTIVE;
assign #(in_delay) CPMC405CPUCLKEN_delay = CPMC405CPUCLKEN;
assign #(in_delay) CPMC405JTAGCLKEN_delay = CPMC405JTAGCLKEN;
assign #(in_delay) CPMC405TIMERCLKEN_delay = CPMC405TIMERCLKEN;
assign #(in_delay) CPMC405TIMERTICK_delay = CPMC405TIMERTICK;
assign #(in_delay) DBGC405DEBUGHALT_delay = DBGC405DEBUGHALT;
assign #(in_delay) DBGC405EXTBUSHOLDACK_delay = DBGC405EXTBUSHOLDACK;
assign #(in_delay) DBGC405UNCONDDEBUGEVENT_delay = DBGC405UNCONDDEBUGEVENT;
assign #(in_delay) DCRC405ACK_delay = DCRC405ACK;
assign #(in_delay) DCRC405DBUSIN_delay[0:31] = DCRC405DBUSIN[0:31];
assign #(in_delay) DSARCVALUE_delay[0:7] = DSARCVALUE[0:7];
assign #(in_delay) DSCNTLVALUE_delay[0:7] = DSCNTLVALUE[0:7];
assign #(in_delay) EICC405CRITINPUTIRQ_delay = EICC405CRITINPUTIRQ;
assign #(in_delay) EICC405EXTINPUTIRQ_delay = EICC405EXTINPUTIRQ;
assign #(in_delay) ISARCVALUE_delay[0:7] = ISARCVALUE[0:7];
assign #(in_delay) ISCNTLVALUE_delay[0:7] = ISCNTLVALUE[0:7];
assign #(in_delay) JTGC405BNDSCANTDO_delay = JTGC405BNDSCANTDO;
assign #(in_delay) JTGC405TCK_delay = JTGC405TCK;
assign #(in_delay) JTGC405TDI_delay = JTGC405TDI;
assign #(in_delay) JTGC405TMS_delay = JTGC405TMS;
assign #(in_delay) JTGC405TRSTNEG_delay = JTGC405TRSTNEG;
assign #(in_delay) MCBCPUCLKEN_delay = MCBCPUCLKEN;
assign #(in_delay) MCBJTAGEN_delay = MCBJTAGEN;
assign #(in_delay) MCBTIMEREN_delay = MCBTIMEREN;
assign #(in_delay) MCPPCRST_delay = MCPPCRST;
assign #(in_delay) PLBC405DCUADDRACK_delay = PLBC405DCUADDRACK;
assign #(in_delay) PLBC405DCUBUSY_delay = PLBC405DCUBUSY;
assign #(in_delay) PLBC405DCUERR_delay = PLBC405DCUERR;
assign #(in_delay) PLBC405DCURDDACK_delay = PLBC405DCURDDACK;
assign #(in_delay) PLBC405DCURDDBUS_delay[0:63] = PLBC405DCURDDBUS[0:63];
assign #(in_delay) PLBC405DCURDWDADDR_delay[1:3] = PLBC405DCURDWDADDR[1:3];
assign #(in_delay) PLBC405DCUSSIZE1_delay = PLBC405DCUSSIZE1;
assign #(in_delay) PLBC405DCUWRDACK_delay = PLBC405DCUWRDACK;
assign #(in_delay) PLBC405ICUADDRACK_delay = PLBC405ICUADDRACK;
assign #(in_delay) PLBC405ICUBUSY_delay = PLBC405ICUBUSY;
assign #(in_delay) PLBC405ICUERR_delay = PLBC405ICUERR;
assign #(in_delay) PLBC405ICURDDACK_delay = PLBC405ICURDDACK;
assign #(in_delay) PLBC405ICURDDBUS_delay[0:63] = PLBC405ICURDDBUS[0:63];
assign #(in_delay) PLBC405ICURDWDADDR_delay[1:3] = PLBC405ICURDWDADDR[1:3];
assign #(in_delay) PLBC405ICUSSIZE1_delay = PLBC405ICUSSIZE1;
assign #(in_delay) RSTC405RESETCHIP_delay = RSTC405RESETCHIP;
assign #(in_delay) RSTC405RESETCORE_delay = RSTC405RESETCORE;
assign #(in_delay) RSTC405RESETSYS_delay = RSTC405RESETSYS;
assign #(in_delay) TIEC405DETERMINISTICMULT_delay = TIEC405DETERMINISTICMULT;
assign #(in_delay) TIEC405DISOPERANDFWD_delay = TIEC405DISOPERANDFWD;
assign #(in_delay) TIEC405MMUEN_delay = TIEC405MMUEN;
assign #(in_delay) TIEDSOCMDCRADDR_delay[0:7] = TIEDSOCMDCRADDR[0:7];
assign #(in_delay) TIEISOCMDCRADDR_delay[0:7] = TIEISOCMDCRADDR[0:7];
assign #(in_delay) TRCC405TRACEDISABLE_delay = TRCC405TRACEDISABLE;
assign #(in_delay) TRCC405TRIGGEREVENTIN_delay = TRCC405TRIGGEREVENTIN;

assign #(out_delay) C405CPMCORESLEEPREQ = C405CPMCORESLEEPREQ_delay;
assign #(out_delay) C405CPMMSRCE = C405CPMMSRCE_delay;
assign #(out_delay) C405CPMMSREE = C405CPMMSREE_delay;
assign #(out_delay) C405CPMTIMERIRQ = C405CPMTIMERIRQ_delay;
assign #(out_delay) C405CPMTIMERRESETREQ = C405CPMTIMERRESETREQ_delay;
assign #(out_delay) C405DBGMSRWE = C405DBGMSRWE_delay;
assign #(out_delay) C405DBGSTOPACK = C405DBGSTOPACK_delay;
assign #(out_delay) C405DBGWBCOMPLETE = C405DBGWBCOMPLETE_delay;
assign #(out_delay) C405DBGWBFULL = C405DBGWBFULL_delay;
assign #(out_delay) C405DBGWBIAR[0:29] = C405DBGWBIAR_delay[0:29];
assign #(out_delay) C405DCRABUS[0:9] = C405DCRABUS_delay[0:9];
assign #(out_delay) C405DCRDBUSOUT[0:31] = C405DCRDBUSOUT_delay[0:31];
assign #(out_delay) C405DCRREAD = C405DCRREAD_delay;
assign #(out_delay) C405DCRWRITE = C405DCRWRITE_delay;
assign #(out_delay) C405JTGCAPTUREDR = C405JTGCAPTUREDR_delay;
assign #(out_delay) C405JTGEXTEST = C405JTGEXTEST_delay;
assign #(out_delay) C405JTGPGMOUT = C405JTGPGMOUT_delay;
assign #(out_delay) C405JTGSHIFTDR = C405JTGSHIFTDR_delay;
assign #(out_delay) C405JTGTDO = C405JTGTDO_delay;
assign #(out_delay) C405JTGTDOEN = C405JTGTDOEN_delay;
assign #(out_delay) C405JTGUPDATEDR = C405JTGUPDATEDR_delay;
assign #(out_delay) C405PLBDCUABORT = C405PLBDCUABORT_delay;
assign #(out_delay) C405PLBDCUABUS[0:31] = C405PLBDCUABUS_delay[0:31];
assign #(out_delay) C405PLBDCUBE[0:7] = C405PLBDCUBE_delay[0:7];
assign #(out_delay) C405PLBDCUCACHEABLE = C405PLBDCUCACHEABLE_delay;
assign #(out_delay) C405PLBDCUGUARDED = C405PLBDCUGUARDED_delay;
assign #(out_delay) C405PLBDCUPRIORITY[0:1] = C405PLBDCUPRIORITY_delay[0:1];
assign #(out_delay) C405PLBDCUREQUEST = C405PLBDCUREQUEST_delay;
assign #(out_delay) C405PLBDCURNW = C405PLBDCURNW_delay;
assign #(out_delay) C405PLBDCUSIZE2 = C405PLBDCUSIZE2_delay;
assign #(out_delay) C405PLBDCUU0ATTR = C405PLBDCUU0ATTR_delay;
assign #(out_delay) C405PLBDCUWRDBUS[0:63] = C405PLBDCUWRDBUS_delay[0:63];
assign #(out_delay) C405PLBDCUWRITETHRU = C405PLBDCUWRITETHRU_delay;
assign #(out_delay) C405PLBICUABORT = C405PLBICUABORT_delay;
assign #(out_delay) C405PLBICUABUS[0:29] = C405PLBICUABUS_delay[0:29];
assign #(out_delay) C405PLBICUCACHEABLE = C405PLBICUCACHEABLE_delay;
assign #(out_delay) C405PLBICUPRIORITY[0:1] = C405PLBICUPRIORITY_delay[0:1];
assign #(out_delay) C405PLBICUREQUEST = C405PLBICUREQUEST_delay;
assign #(out_delay) C405PLBICUSIZE[2:3] = C405PLBICUSIZE_delay[2:3];
assign #(out_delay) C405PLBICUU0ATTR = C405PLBICUU0ATTR_delay;
assign #(out_delay) C405RSTCHIPRESETREQ = C405RSTCHIPRESETREQ_delay;
assign #(out_delay) C405RSTCORERESETREQ = C405RSTCORERESETREQ_delay;
assign #(out_delay) C405RSTSYSRESETREQ = C405RSTSYSRESETREQ_delay;
assign #(out_delay) C405TRCCYCLE = C405TRCCYCLE_delay;
assign #(out_delay) C405TRCEVENEXECUTIONSTATUS[0:1] = C405TRCEVENEXECUTIONSTATUS_delay[0:1];
assign #(out_delay) C405TRCODDEXECUTIONSTATUS[0:1] = C405TRCODDEXECUTIONSTATUS_delay[0:1];
assign #(out_delay) C405TRCTRACESTATUS[0:3] = C405TRCTRACESTATUS_delay[0:3];
assign #(out_delay) C405TRCTRIGGEREVENTOUT = C405TRCTRIGGEREVENTOUT_delay;
assign #(out_delay) C405TRCTRIGGEREVENTTYPE[0:10] = C405TRCTRIGGEREVENTTYPE_delay[0:10];
assign #(out_delay) C405XXXMACHINECHECK = C405XXXMACHINECHECK_delay;
assign #(out_delay) DSOCMBRAMABUS[8:29] = DSOCMBRAMABUS_delay[8:29];
assign #(out_delay) DSOCMBRAMBYTEWRITE[0:3] = DSOCMBRAMBYTEWRITE_delay[0:3];
assign #(out_delay) DSOCMBRAMEN = DSOCMBRAMEN_delay;
assign #(out_delay) DSOCMBRAMWRDBUS[0:31] = DSOCMBRAMWRDBUS_delay[0:31];
assign #(out_delay) DSOCMBUSY = DSOCMBUSY_delay;
assign #(out_delay) ISOCMBRAMEN = ISOCMBRAMEN_delay;
assign #(out_delay) ISOCMBRAMEVENWRITEEN = ISOCMBRAMEVENWRITEEN_delay;
assign #(out_delay) ISOCMBRAMODDWRITEEN = ISOCMBRAMODDWRITEEN_delay;
assign #(out_delay) ISOCMBRAMRDABUS[8:28] = ISOCMBRAMRDABUS_delay[8:28];
assign #(out_delay) ISOCMBRAMWRABUS[8:28] = ISOCMBRAMWRABUS_delay[8:28];
assign #(out_delay) ISOCMBRAMWRDBUS[0:31] = ISOCMBRAMWRDBUS_delay[0:31];

wire    FPGA_CCLK;
wire	FPGA_BUS_RESET;
wire	FPGA_GSR;
wire	FPGA_GWE;
wire	FPGA_GHIGHB;
wire	GSR_OR;

reg	FPGA_POR;
reg	FPGA_CCLK_REG;

tri0 GSR = glbl.GSR;

`ifdef STARTUP_BLK
	assign FPGA_CCLK	= TESTBENCH.FPGA_cclk;
	assign  FPGA_BUS_RESET 	= TESTBENCH.FPGA_bus_reset;
	assign  GSR_OR 		= TESTBENCH.FPGA_gsr;
	assign  FPGA_GWE 	= TESTBENCH.FPGA_gwe;
	assign  FPGA_GHIGHB 	= TESTBENCH.FPGA_ghigh_b;
`else

FPGA_startup start_blk(
.bus_reset	(FPGA_BUS_RESET),
.ghigh_b	(FPGA_GHIGHB), 
.gsr		(FPGA_GSR), 
.done		(), 
.gwe		(FPGA_GWE), 
.gts_b		(), 
.shutdown	(1'b0), 
.cclk		(FPGA_CCLK), 
.por		(FPGA_POR)
);

or IGSR_OR (GSR_OR, FPGA_GSR, GSR);

`define Loc_FPGA_POR_TIME           100   // FPGA Power-On Reset time

// Generate FPGA CCLK
 always
    #5000 FPGA_CCLK_REG = ~FPGA_CCLK_REG;

assign FPGA_CCLK = FPGA_CCLK_REG;

initial begin
    FPGA_CCLK_REG = 0;
    FPGA_POR  = 1'b1;
    #(`Loc_FPGA_POR_TIME)       FPGA_POR  = 1'b0;
end

`endif   // STARTUP_BLK

wire FPGA_BUS_RESET_delay;
wire GSR_delay;
wire FPGA_GWE_delay;
wire FPGA_GHIGHB_delay;

assign #(in_delay) FPGA_BUS_RESET_delay = FPGA_BUS_RESET;
assign #(in_delay) GSR_delay = GSR_OR;
assign #(in_delay) FPGA_GWE_delay = FPGA_GWE;
assign #(in_delay) FPGA_GHIGHB_delay = FPGA_GHIGHB;

`ifdef ProcBlk_RTL
usr_proc_block_cap Iusr_proc_block_cap(
`else
PPC405_SWIFT IPPC405_SWIFT(
`endif          //ProcBlk_rtl

   .BUS_CLK(FPGA_CCLK),
   .BUS_RESET(FPGA_BUS_RESET_delay),
   .GSR(GSR_delay),
   .GWE(FPGA_GWE_delay),
   .GHIGHB(FPGA_GHIGHB_delay),
   .CPMC405CPUCLKEN(CPMC405CPUCLKEN_delay),
   .CPMC405JTAGCLKEN(CPMC405JTAGCLKEN_delay),
   .CPMC405TIMERCLKEN(CPMC405TIMERCLKEN_delay),
   .C405JTGPGMOUT(C405JTGPGMOUT_delay),
   .MCBCPUCLKEN(MCBCPUCLKEN_delay),
   .MCBJTAGEN(MCBJTAGEN_delay),
   .MCBTIMEREN(MCBTIMEREN_delay),
   .MCPPCRST(MCPPCRST_delay),
   .C405TRCODDEXECUTIONSTATUS(C405TRCODDEXECUTIONSTATUS_delay),
   .C405TRCEVENEXECUTIONSTATUS(C405TRCEVENEXECUTIONSTATUS_delay),
   .CPMC405CLOCK(CPMC405CLOCK),
   .CPMC405CORECLKINACTIVE(CPMC405CORECLKINACTIVE_delay),
   .PLBCLK(PLBCLK),
   .CPMC405TIMERTICK(CPMC405TIMERTICK_delay),
   .C405CPMMSREE(C405CPMMSREE_delay),
   .C405CPMMSRCE(C405CPMMSRCE_delay),
   .C405CPMTIMERIRQ(C405CPMTIMERIRQ_delay),
   .C405CPMTIMERRESETREQ(C405CPMTIMERRESETREQ_delay),
   .C405CPMCORESLEEPREQ(C405CPMCORESLEEPREQ_delay),
   .TIEC405DISOPERANDFWD(TIEC405DISOPERANDFWD_delay),
   .TIEC405DETERMINISTICMULT(TIEC405DETERMINISTICMULT_delay),
   .TIEC405MMUEN(TIEC405MMUEN_delay),
   .TIEC405PVR(PPCUSER),
   .C405XXXMACHINECHECK(C405XXXMACHINECHECK_delay),
   .C405RSTCHIPRESETREQ(C405RSTCHIPRESETREQ_delay),
   .C405RSTCORERESETREQ(C405RSTCORERESETREQ_delay),
   .C405RSTSYSRESETREQ(C405RSTSYSRESETREQ_delay),
   .RSTC405RESETCHIP(RSTC405RESETCHIP_delay),
   .RSTC405RESETCORE(RSTC405RESETCORE_delay),
   .RSTC405RESETSYS(RSTC405RESETSYS_delay),
   .C405PLBICUREQUEST(C405PLBICUREQUEST_delay),
   .C405PLBICUPRIORITY(C405PLBICUPRIORITY_delay),
   .C405PLBICUCACHEABLE(C405PLBICUCACHEABLE_delay),
   .C405PLBICUABUS(C405PLBICUABUS_delay),
   .C405PLBICUSIZE(C405PLBICUSIZE_delay),
   .C405PLBICUABORT(C405PLBICUABORT_delay),
   .C405PLBICUU0ATTR(C405PLBICUU0ATTR_delay),
   .PLBC405ICUADDRACK(PLBC405ICUADDRACK_delay),
   .PLBC405ICUBUSY(PLBC405ICUBUSY_delay),
   .PLBC405ICUERR(PLBC405ICUERR_delay),
   .PLBC405ICURDDACK(PLBC405ICURDDACK_delay),
   .PLBC405ICURDDBUS(PLBC405ICURDDBUS_delay),
   .PLBC405ICUSSIZE1(PLBC405ICUSSIZE1_delay),
   .PLBC405ICURDWDADDR(PLBC405ICURDWDADDR_delay),
   .C405PLBDCUREQUEST(C405PLBDCUREQUEST_delay),
   .C405PLBDCURNW(C405PLBDCURNW_delay),
   .C405PLBDCUABUS(C405PLBDCUABUS_delay),
   .C405PLBDCUBE(C405PLBDCUBE_delay),
   .C405PLBDCUCACHEABLE(C405PLBDCUCACHEABLE_delay),
   .C405PLBDCUGUARDED(C405PLBDCUGUARDED_delay),
   .C405PLBDCUPRIORITY(C405PLBDCUPRIORITY_delay),
   .C405PLBDCUSIZE2(C405PLBDCUSIZE2_delay),
   .C405PLBDCUABORT(C405PLBDCUABORT_delay),
   .C405PLBDCUWRDBUS(C405PLBDCUWRDBUS_delay),
   .C405PLBDCUU0ATTR(C405PLBDCUU0ATTR_delay),
   .C405PLBDCUWRITETHRU(C405PLBDCUWRITETHRU_delay),
   .PLBC405DCUADDRACK(PLBC405DCUADDRACK_delay),
   .PLBC405DCUBUSY(PLBC405DCUBUSY_delay),
   .PLBC405DCUERR(PLBC405DCUERR_delay),
   .PLBC405DCURDDACK(PLBC405DCURDDACK_delay),
   .PLBC405DCURDDBUS(PLBC405DCURDDBUS_delay),
   .PLBC405DCURDWDADDR(PLBC405DCURDWDADDR_delay),
   .PLBC405DCUSSIZE1(PLBC405DCUSSIZE1_delay),
   .PLBC405DCUWRDACK(PLBC405DCUWRDACK_delay),
   .ISOCMBRAMRDABUS(ISOCMBRAMRDABUS_delay),
   .ISOCMBRAMWRABUS(ISOCMBRAMWRABUS_delay),
   .ISOCMBRAMEN(ISOCMBRAMEN_delay),
   .ISOCMBRAMODDWRITEEN(ISOCMBRAMODDWRITEEN_delay),
   .ISOCMBRAMEVENWRITEEN(ISOCMBRAMEVENWRITEEN_delay),
   .ISOCMBRAMWRDBUS(ISOCMBRAMWRDBUS_delay),
   .BRAMISOCMRDDBUS(BRAMISOCMRDDBUS_delay),
   .TIEISOCMDCRADDR(TIEISOCMDCRADDR_delay),
   .ISARCVALUE(ISARCVALUE_delay),
   .ISCNTLVALUE(ISCNTLVALUE_delay),
   .BRAMISOCMCLK(BRAMISOCMCLK),
   .DSOCMBRAMABUS(DSOCMBRAMABUS_delay),
   .DSOCMBRAMBYTEWRITE(DSOCMBRAMBYTEWRITE_delay),
   .DSOCMBRAMEN(DSOCMBRAMEN_delay),
   .DSOCMBRAMWRDBUS(DSOCMBRAMWRDBUS_delay),
   .BRAMDSOCMRDDBUS(BRAMDSOCMRDDBUS_delay),
   .DSOCMBUSY(DSOCMBUSY_delay),
   .TIEDSOCMDCRADDR(TIEDSOCMDCRADDR_delay),
   .DSARCVALUE(DSARCVALUE_delay),
   .DSCNTLVALUE(DSCNTLVALUE_delay),
   .BRAMDSOCMCLK(BRAMDSOCMCLK),
   .C405DCRREAD(C405DCRREAD_delay),
   .C405DCRWRITE(C405DCRWRITE_delay),
   .C405DCRABUS(C405DCRABUS_delay),
   .C405DCRDBUSOUT(C405DCRDBUSOUT_delay),
   .DCRC405ACK(DCRC405ACK_delay),
   .DCRC405DBUSIN(DCRC405DBUSIN_delay),
   .EICC405EXTINPUTIRQ(EICC405EXTINPUTIRQ_delay),
   .EICC405CRITINPUTIRQ(EICC405CRITINPUTIRQ_delay),
   .JTGC405BNDSCANTDO(JTGC405BNDSCANTDO_delay),
   .JTGC405TCK(JTGC405TCK_delay),
   .JTGC405TDI(JTGC405TDI_delay),
   .JTGC405TMS(JTGC405TMS_delay),
   .JTGC405TRSTNEG(JTGC405TRSTNEG_delay),
   .C405JTGTDO(C405JTGTDO_delay),
   .C405JTGTDOEN(C405JTGTDOEN_delay),
   .C405JTGEXTEST(C405JTGEXTEST_delay),
   .C405JTGCAPTUREDR(C405JTGCAPTUREDR_delay),
   .C405JTGSHIFTDR(C405JTGSHIFTDR_delay),
   .C405JTGUPDATEDR(C405JTGUPDATEDR_delay),
   .DBGC405DEBUGHALT(DBGC405DEBUGHALT_delay),
   .DBGC405UNCONDDEBUGEVENT(DBGC405UNCONDDEBUGEVENT_delay),
   .DBGC405EXTBUSHOLDACK(DBGC405EXTBUSHOLDACK_delay),
   .C405DBGMSRWE(C405DBGMSRWE_delay),
   .C405DBGSTOPACK(C405DBGSTOPACK_delay),
   .C405DBGWBCOMPLETE(C405DBGWBCOMPLETE_delay),
   .C405DBGWBFULL(C405DBGWBFULL_delay),
   .C405DBGWBIAR(C405DBGWBIAR_delay),
   .C405TRCTRIGGEREVENTOUT(C405TRCTRIGGEREVENTOUT_delay),
   .C405TRCTRIGGEREVENTTYPE(C405TRCTRIGGEREVENTTYPE_delay),
   .C405TRCCYCLE(C405TRCCYCLE_delay),
   .C405TRCTRACESTATUS(C405TRCTRACESTATUS_delay),
   .TRCC405TRACEDISABLE(TRCC405TRACEDISABLE_delay),
   .TRCC405TRIGGEREVENTIN(TRCC405TRIGGEREVENTIN_delay)
);

endmodule

module FPGA_startup(bus_reset, ghigh_b, gsr, done, gwe, gts_b, shutdown, cclk, por);
   output bus_reset;
   output ghigh_b;
   output gsr;
   output done;
   output gwe;
   output gts_b;
   input  shutdown;
   input  cclk, por;

   reg    bus_reset, abus_reset;
   reg    ghigh_b, aghigh_b;
   reg    gsr, agsr;
   reg    done, adone;
   reg    gwe, agwe;
   reg    gts_b, agts_b;

   reg    [7:0] count;

   always @ (posedge cclk or posedge por) begin
     if(por) count <= {8{1'b0}};
     else if(shutdown && (count > {8{1'b0}})) count = count - 1;
     else if(!shutdown && (count < {8'hFF})) count = count + 1;
   end

   always @ (posedge cclk or posedge por) begin
     if(por) begin
       {bus_reset,ghigh_b,gsr,done,gwe,gts_b} <= 6'b100000;
     end else begin
       {bus_reset,ghigh_b,gsr,done,gwe,gts_b} <= 
                                   {abus_reset,aghigh_b,agsr,adone,agwe,agts_b};
     end
   end

   always @ (count) begin
     // defaults
     
     abus_reset = 1;
     aghigh_b = 0;
     agsr = 0;
     adone = 0;
     agwe = 0;
     agts_b = 0;

     // Trip times are in order for default sequence.
     if(count >= 8'h04) abus_reset = 0;
     if(count == 8'h21 || count == 8'h22) agsr = 1;
     if(count > 8'h26) aghigh_b = 1;
     if(count > 8'h31) adone = 1;
     if(count > 8'h32) agwe = 1;
     if(count > 8'h33) agts_b = 1;
   end
   
endmodule // startup
