
/*

FUNCTION	: VCC cell

*/

`timescale  100 ps / 10 ps

`celldefine

module VCC(P);


    output P;

	assign P = 1'b1;

endmodule

`endcelldefine
