// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CAPTURE_FPGACORE.v,v 1.1 2003/01/23 01:39:09 wloo Exp $
/*

FUNCTION	: Special Function Cell, CAPTURE_FPGACORE

*/

`timescale  100 ps / 10 ps


module CAPTURE_FPGACORE (CAP, CLK);

    input  CAP, CLK;

endmodule

