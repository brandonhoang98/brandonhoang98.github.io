//    Xilinx Proprietary Primitive Cell X_ZERO for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_ZERO.v,v 1.10 2003/01/21 02:38:45 wloo Exp $
//

`timescale 1 ps/1 ps

module X_ZERO (O);

  output O;

  assign O = 1'b0;

endmodule
