// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/TBLOCK.v,v 1.8 2003/01/21 01:55:44 wloo Exp $

/*

FUNCTION	: TBLOCK dummy simulation module

*/

`timescale  100 ps / 10 ps


module TBLOCK ();

endmodule

