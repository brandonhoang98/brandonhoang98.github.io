// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CAPTURE_SPARTAN3.v,v 1.2 2003/01/21 01:55:23 wloo Exp $
/*

FUNCTION	: Special Function Cell, CAPTURE_SPARTAN3

*/

`timescale  100 ps / 10 ps


module CAPTURE_SPARTAN3 (CAP, CLK);

    input  CAP, CLK;

endmodule

