
/*

FUNCTION	: TIMEGRP dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module TIMEGRP ();


endmodule

`endcelldefine
