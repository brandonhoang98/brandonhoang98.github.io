//    Xilinx Proprietary Primitive Cell X_XOR32 for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_XOR32.v,v 1.9 2003/01/21 02:38:45 wloo Exp $
//

`timescale 1 ps/1 ps

module X_XOR32 (O, I0, I1, I2, I3, I4, I5, I6, I7,
                I8, I9, I10, I11, I12, I13, I14, I15,
                I16, I17, I18, I19, I20, I21, I22, I23,
                I24, I25, I26, I27, I28, I29, I30, I31);

  output O;
  input I0, I1, I2, I3, I4, I5, I6, I7,
        I8, I9, I10, I11, I12, I13, I14, I15,
        I16, I17, I18, I19, I20, I21, I22, I23,
        I24, I25, I26, I27, I28, I29, I30, I31;

  xor (O, I0, I1, I2, I3, I4, I5, I6, I7,
       I8, I9, I10, I11, I12, I13, I14, I15,
       I16, I17, I18, I19, I20, I21, I22, I23,
       I24, I25, I26, I27, I28, I29, I30, I31);

  specify

	(I0 => O) = (0:0:0, 0:0:0);
	(I1 => O) = (0:0:0, 0:0:0);
	(I2 => O) = (0:0:0, 0:0:0);
	(I3 => O) = (0:0:0, 0:0:0);
	(I4 => O) = (0:0:0, 0:0:0);
	(I5 => O) = (0:0:0, 0:0:0);
	(I6 => O) = (0:0:0, 0:0:0);
	(I7 => O) = (0:0:0, 0:0:0);
	(I8 => O) = (0:0:0, 0:0:0);
	(I9 => O) = (0:0:0, 0:0:0);
	(I10 => O) = (0:0:0, 0:0:0);
	(I11 => O) = (0:0:0, 0:0:0);
	(I12 => O) = (0:0:0, 0:0:0);
	(I13 => O) = (0:0:0, 0:0:0);
	(I14 => O) = (0:0:0, 0:0:0);
	(I15 => O) = (0:0:0, 0:0:0);
	(I16 => O) = (0:0:0, 0:0:0);
	(I17 => O) = (0:0:0, 0:0:0);
	(I18 => O) = (0:0:0, 0:0:0);
	(I19 => O) = (0:0:0, 0:0:0);
	(I20 => O) = (0:0:0, 0:0:0);
	(I21 => O) = (0:0:0, 0:0:0);
	(I22 => O) = (0:0:0, 0:0:0);
	(I23 => O) = (0:0:0, 0:0:0);
	(I24 => O) = (0:0:0, 0:0:0);
	(I25 => O) = (0:0:0, 0:0:0);
	(I26 => O) = (0:0:0, 0:0:0);
	(I27 => O) = (0:0:0, 0:0:0);
	(I28 => O) = (0:0:0, 0:0:0);
	(I29 => O) = (0:0:0, 0:0:0);
	(I30 => O) = (0:0:0, 0:0:0);
	(I31 => O) = (0:0:0, 0:0:0);

	specparam PATHPULSE$ = 0;

  endspecify

endmodule
