
/*

FUNCTION	: TIMESPEC dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module TIMESPEC ();


endmodule

`endcelldefine
