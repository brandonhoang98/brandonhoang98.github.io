//    Xilinx Proprietary Primitive Cell X_BPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_BPAD.v,v 1.9 2003/01/21 02:38:33 wloo Exp $
//

`timescale 1 ps/1 ps

module X_BPAD (PAD);

  inout PAD;

endmodule
