//    Xilinx Proprietary Primitive Cell X_ONE for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_ONE.v,v 1.10 2003/01/21 02:38:37 wloo Exp $
//

`timescale 1 ps/1 ps

module X_ONE (O);

  output O;

  assign O = 1'b1;

endmodule
