
/*

FUNCTION	: TBLOCK dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module TBLOCK ();


endmodule

`endcelldefine
