//    Xilinx Proprietary Primitive Cell X_IPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_IPAD.v,v 1.9 2003/01/21 02:38:36 wloo Exp $
//

`timescale 1 ps/1 ps

module X_IPAD (PAD);

  input PAD;

endmodule
