
/*

FUNCTION	: MERGE dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module MERGE (I);


    input  I;

endmodule

`endcelldefine
