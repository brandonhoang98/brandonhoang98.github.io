
/*

FUNCTION	: MIN_OFF dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module MIN_OFF (I);


    input  I;

endmodule

`endcelldefine
