// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/GND.v,v 1.8 2003/01/21 01:55:23 wloo Exp $

/*

FUNCTION	: GND cell

*/

`timescale  100 ps / 10 ps


module GND(G);

    output G;

	assign G = 1'b0;

endmodule

