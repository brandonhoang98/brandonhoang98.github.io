
/*

FUNCTION	: OPT_UIM dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module OPT_UIM (I);


    input  I;

endmodule

`endcelldefine
