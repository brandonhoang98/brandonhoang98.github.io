
/*

FUNCTION	: KEEP dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module KEEP (O, I);


    output O;

    input  I;

endmodule

`endcelldefine
