//    Xilinx Proprietary Primitive Cell X_OPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_OPAD.v,v 1.9 2003/01/21 02:38:37 wloo Exp $
//

`timescale 1 ps/1 ps

module X_OPAD (PAD);

  output PAD;

endmodule
