// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/CONFIG.v,v 1.8 2003/01/21 01:55:23 wloo Exp $

/*

FUNCTION	: CONFIG dummy simulation module

*/

`timescale  100 ps / 10 ps


module CONFIG ();

endmodule

