
/*

FUNCTION	: WIREAND dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module WIREAND (I);


    input  I;

endmodule

`endcelldefine
