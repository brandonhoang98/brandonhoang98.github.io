// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/verunilibs/s/FMAP.v,v 1.8 2003/01/21 01:55:23 wloo Exp $

/*

FUNCTION	: FMAP dummy simulation module

*/

`timescale  100 ps / 10 ps


module FMAP (I1, I2, I3, I4, O);

    input  I1, I2, I3, I4, O;

endmodule

