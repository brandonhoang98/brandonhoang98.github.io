
/*

FUNCTION	: GND cell

*/

`timescale  100 ps / 10 ps

`celldefine

module GND(G);


    output G;

	assign G = 1'b0;

endmodule

`endcelldefine
