// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_PPC405.v,v 1.15 2003/01/21 02:38:38 wloo Exp $

/*

		: Power PC

*/

`timescale  1 ps / 1 ps

module X_PPC405 (
		C405CPMCORESLEEPREQ,
		C405CPMMSRCE,
		C405CPMMSREE,
		C405CPMTIMERIRQ,
		C405CPMTIMERRESETREQ,
		C405DBGMSRWE,
		C405DBGSTOPACK,
		C405DBGWBCOMPLETE,
		C405DBGWBFULL,
		C405DBGWBIAR,
		C405DCRABUS,
		C405DCRDBUSOUT,
		C405DCRREAD,
		C405DCRWRITE,
		C405JTGCAPTUREDR,
		C405JTGEXTEST,
		C405JTGPGMOUT,
		C405JTGSHIFTDR,
		C405JTGTDO,
		C405JTGTDOEN,
		C405JTGUPDATEDR,
		C405PLBDCUABORT,
		C405PLBDCUABUS,
		C405PLBDCUBE,
		C405PLBDCUCACHEABLE,
		C405PLBDCUGUARDED,
		C405PLBDCUPRIORITY,
		C405PLBDCUREQUEST,
		C405PLBDCURNW,
		C405PLBDCUSIZE2,
		C405PLBDCUU0ATTR,
		C405PLBDCUWRDBUS,
		C405PLBDCUWRITETHRU,
		C405PLBICUABORT,
		C405PLBICUABUS,
		C405PLBICUCACHEABLE,
		C405PLBICUPRIORITY,
		C405PLBICUREQUEST,
		C405PLBICUSIZE,
		C405PLBICUU0ATTR,
		C405RSTCHIPRESETREQ,
		C405RSTCORERESETREQ,
		C405RSTSYSRESETREQ,
		C405TRCCYCLE,
		C405TRCEVENEXECUTIONSTATUS,
		C405TRCODDEXECUTIONSTATUS,
		C405TRCTRACESTATUS,
		C405TRCTRIGGEREVENTOUT,
		C405TRCTRIGGEREVENTTYPE,
		C405XXXMACHINECHECK,
		DSOCMBRAMABUS,
		DSOCMBRAMBYTEWRITE,
		DSOCMBRAMEN,
		DSOCMBRAMWRDBUS,
		DSOCMBUSY,
		ISOCMBRAMEN,
		ISOCMBRAMEVENWRITEEN,
		ISOCMBRAMODDWRITEEN,
		ISOCMBRAMRDABUS,
		ISOCMBRAMWRABUS,
		ISOCMBRAMWRDBUS,

		BRAMDSOCMCLK,
		BRAMDSOCMRDDBUS,
		BRAMISOCMCLK,
		BRAMISOCMRDDBUS,
		CPMC405CLOCK,
		CPMC405CORECLKINACTIVE,
		CPMC405CPUCLKEN,
		CPMC405JTAGCLKEN,
		CPMC405TIMERCLKEN,
		CPMC405TIMERTICK,
		DBGC405DEBUGHALT,
		DBGC405EXTBUSHOLDACK,
		DBGC405UNCONDDEBUGEVENT,
		DCRC405ACK,
		DCRC405DBUSIN,
		DSARCVALUE,
		DSCNTLVALUE,
		EICC405CRITINPUTIRQ,
		EICC405EXTINPUTIRQ,
		GSR,
		ISARCVALUE,
		ISCNTLVALUE,
		JTGC405BNDSCANTDO,
		JTGC405TCK,
		JTGC405TDI,
		JTGC405TMS,
		JTGC405TRSTNEG,
		MCBCPUCLKEN,
		MCBJTAGEN,
		MCBTIMEREN,
		MCPPCRST,
		PLBC405DCUADDRACK,
		PLBC405DCUBUSY,
		PLBC405DCUERR,
		PLBC405DCURDDACK,
		PLBC405DCURDDBUS,
		PLBC405DCURDWDADDR,
		PLBC405DCUSSIZE1,
		PLBC405DCUWRDACK,
		PLBC405ICUADDRACK,
		PLBC405ICUBUSY,
		PLBC405ICUERR,
		PLBC405ICURDDACK,
		PLBC405ICURDDBUS,
		PLBC405ICURDWDADDR,
		PLBC405ICUSSIZE1,
		PLBCLK,
		RSTC405RESETCHIP,
		RSTC405RESETCORE,
		RSTC405RESETSYS,
		TIEC405DETERMINISTICMULT,
		TIEC405DISOPERANDFWD,
		TIEC405MMUEN,
		TIEDSOCMDCRADDR,
		TIEISOCMDCRADDR,
		TRCC405TRACEDISABLE,
		TRCC405TRIGGEREVENTIN
);

parameter in_delay=0;
parameter out_delay=0;
parameter PPCUSER = 4'b0000;

output		C405CPMCORESLEEPREQ;
output		C405CPMMSRCE;
output		C405CPMMSREE;
output		C405CPMTIMERIRQ;
output		C405CPMTIMERRESETREQ;
output		C405DBGMSRWE;
output		C405DBGSTOPACK;
output		C405DBGWBCOMPLETE;
output		C405DBGWBFULL;
output	[0:29]	C405DBGWBIAR;
output	[0:9]	C405DCRABUS;
output	[0:31]	C405DCRDBUSOUT;
output		C405DCRREAD;
output		C405DCRWRITE;
output		C405JTGCAPTUREDR;
output		C405JTGEXTEST;
output		C405JTGPGMOUT;
output		C405JTGSHIFTDR;
output		C405JTGTDO;
output		C405JTGTDOEN;
output		C405JTGUPDATEDR;
output		C405PLBDCUABORT;
output	[0:31]	C405PLBDCUABUS;
output	[0:7]	C405PLBDCUBE;
output		C405PLBDCUCACHEABLE;
output		C405PLBDCUGUARDED;
output	[0:1]	C405PLBDCUPRIORITY;
output		C405PLBDCUREQUEST;
output		C405PLBDCURNW;
output		C405PLBDCUSIZE2;
output		C405PLBDCUU0ATTR;
output	[0:63]	C405PLBDCUWRDBUS;
output		C405PLBDCUWRITETHRU;
output		C405PLBICUABORT;
output	[0:29]	C405PLBICUABUS;
output		C405PLBICUCACHEABLE;
output	[0:1]	C405PLBICUPRIORITY;
output		C405PLBICUREQUEST;
output	[2:3]	C405PLBICUSIZE;
output		C405PLBICUU0ATTR;
output		C405RSTCHIPRESETREQ;
output		C405RSTCORERESETREQ;
output		C405RSTSYSRESETREQ;
output		C405TRCCYCLE;
output	[0:1]	C405TRCEVENEXECUTIONSTATUS;
output	[0:1]	C405TRCODDEXECUTIONSTATUS;
output	[0:3]	C405TRCTRACESTATUS;
output		C405TRCTRIGGEREVENTOUT;
output	[0:10]	C405TRCTRIGGEREVENTTYPE;
output		C405XXXMACHINECHECK;
output	[8:29]	DSOCMBRAMABUS;
output	[0:3]	DSOCMBRAMBYTEWRITE;
output		DSOCMBRAMEN;
output	[0:31]	DSOCMBRAMWRDBUS;
output		DSOCMBUSY;
output		ISOCMBRAMEN;
output		ISOCMBRAMEVENWRITEEN;
output		ISOCMBRAMODDWRITEEN;
output	[8:28]	ISOCMBRAMRDABUS;
output	[8:28]	ISOCMBRAMWRABUS;
output	[0:31]	ISOCMBRAMWRDBUS;

input		BRAMDSOCMCLK;
input	[0:31]	BRAMDSOCMRDDBUS;
input		BRAMISOCMCLK;
input	[0:63]	BRAMISOCMRDDBUS;
input		CPMC405CLOCK;
input		CPMC405CORECLKINACTIVE;
input		CPMC405CPUCLKEN;
input		CPMC405JTAGCLKEN;
input		CPMC405TIMERCLKEN;
input		CPMC405TIMERTICK;
input		DBGC405DEBUGHALT;
input		DBGC405EXTBUSHOLDACK;
input		DBGC405UNCONDDEBUGEVENT;
input		DCRC405ACK;
input	[0:31]	DCRC405DBUSIN;
input	[0:7]	DSARCVALUE;
input	[0:7]	DSCNTLVALUE;
input		EICC405CRITINPUTIRQ;
input		EICC405EXTINPUTIRQ;
input		GSR;
input	[0:7]	ISARCVALUE;
input	[0:7]	ISCNTLVALUE;
input		JTGC405BNDSCANTDO;
input		JTGC405TCK;
input		JTGC405TDI;
input		JTGC405TMS;
input		JTGC405TRSTNEG;
input		MCBCPUCLKEN;
input		MCBJTAGEN;
input		MCBTIMEREN;
input		MCPPCRST;
input		PLBC405DCUADDRACK;
input		PLBC405DCUBUSY;
input		PLBC405DCUERR;
input		PLBC405DCURDDACK;
input	[0:63]	PLBC405DCURDDBUS;
input	[1:3]	PLBC405DCURDWDADDR;
input		PLBC405DCUSSIZE1;
input		PLBC405DCUWRDACK;
input		PLBC405ICUADDRACK;
input		PLBC405ICUBUSY;
input		PLBC405ICUERR;
input		PLBC405ICURDDACK;
input	[0:63]	PLBC405ICURDDBUS;
input	[1:3]	PLBC405ICURDWDADDR;
input		PLBC405ICUSSIZE1;
input		PLBCLK;
input		RSTC405RESETCHIP;
input		RSTC405RESETCORE;
input		RSTC405RESETSYS;
input		TIEC405DETERMINISTICMULT;
input		TIEC405DISOPERANDFWD;
input		TIEC405MMUEN;
input	[0:7]	TIEDSOCMDCRADDR;
input	[0:7]	TIEISOCMDCRADDR;
input		TRCC405TRACEDISABLE;
input		TRCC405TRIGGEREVENTIN;

reg notifier;

// define input delay bus

wire [0:31] BRAMDSOCMRDDBUS_delay;
wire [0:63] BRAMISOCMRDDBUS_delay;
wire [0:31] DCRC405DBUSIN_delay;
wire [0:7] DSARCVALUE_delay;
wire [0:7] DSCNTLVALUE_delay;
wire [0:7] ISARCVALUE_delay;
wire [0:7] ISCNTLVALUE_delay;
wire [0:63] PLBC405DCURDDBUS_delay;
wire [1:3] PLBC405DCURDWDADDR_delay;
wire [0:63] PLBC405ICURDDBUS_delay;
wire [1:3] PLBC405ICURDWDADDR_delay;
wire [0:7] TIEDSOCMDCRADDR_delay;
wire [0:7] TIEISOCMDCRADDR_delay;

// define input delay pins

wire CPMC405CORECLKINACTIVE_delay;
wire CPMC405CPUCLKEN_delay;
wire CPMC405JTAGCLKEN_delay;
wire CPMC405TIMERCLKEN_delay;
wire CPMC405TIMERTICK_delay;
wire DBGC405DEBUGHALT_delay;
wire DBGC405EXTBUSHOLDACK_delay;
wire DBGC405UNCONDDEBUGEVENT_delay;
wire DCRC405ACK_delay;
wire EICC405CRITINPUTIRQ_delay;
wire EICC405EXTINPUTIRQ_delay;
wire JTGC405BNDSCANTDO_delay;
wire JTGC405TCK_delay;
wire JTGC405TDI_delay;
wire JTGC405TMS_delay;
wire JTGC405TRSTNEG_delay;
wire MCBCPUCLKEN_delay;
wire MCBJTAGEN_delay;
wire MCBTIMEREN_delay;
wire MCPPCRST_delay;
wire PLBC405DCUADDRACK_delay;
wire PLBC405DCUBUSY_delay;
wire PLBC405DCUERR_delay;
wire PLBC405DCURDDACK_delay;
wire PLBC405DCUSSIZE1_delay;
wire PLBC405DCUWRDACK_delay;
wire PLBC405ICUADDRACK_delay;
wire PLBC405ICUBUSY_delay;
wire PLBC405ICUERR_delay;
wire PLBC405ICURDDACK_delay;
wire PLBC405ICUSSIZE1_delay;
wire RSTC405RESETCHIP_delay;
wire RSTC405RESETCORE_delay;
wire RSTC405RESETSYS_delay;
wire TIEC405DETERMINISTICMULT_delay;
wire TIEC405DISOPERANDFWD_delay;
wire TIEC405MMUEN_delay;
wire TRCC405TRACEDISABLE_delay;
wire TRCC405TRIGGEREVENTIN_delay;

// define output delay bus

wire [0:29] C405DBGWBIAR_delay;
wire [0:9] C405DCRABUS_delay;
wire [0:31] C405DCRDBUSOUT_delay;
wire [0:31] C405PLBDCUABUS_delay;
wire [0:7] C405PLBDCUBE_delay;
wire [0:1] C405PLBDCUPRIORITY_delay;
wire [0:63] C405PLBDCUWRDBUS_delay;
wire [0:29] C405PLBICUABUS_delay;
wire [0:1] C405PLBICUPRIORITY_delay;
wire [2:3] C405PLBICUSIZE_delay;
wire [0:1] C405TRCEVENEXECUTIONSTATUS_delay;
wire [0:1] C405TRCODDEXECUTIONSTATUS_delay;
wire [0:3] C405TRCTRACESTATUS_delay;
wire [0:10] C405TRCTRIGGEREVENTTYPE_delay;
wire [8:29] DSOCMBRAMABUS_delay;
wire [0:3] DSOCMBRAMBYTEWRITE_delay;
wire [0:31] DSOCMBRAMWRDBUS_delay;
wire [8:28] ISOCMBRAMRDABUS_delay;
wire [8:28] ISOCMBRAMWRABUS_delay;
wire [0:31] ISOCMBRAMWRDBUS_delay;

// define output delay pins

wire C405CPMCORESLEEPREQ_delay;
wire C405CPMMSRCE_delay;
wire C405CPMMSREE_delay;
wire C405CPMTIMERIRQ_delay;
wire C405CPMTIMERRESETREQ_delay;
wire C405DBGMSRWE_delay;
wire C405DBGSTOPACK_delay;
wire C405DBGWBCOMPLETE_delay;
wire C405DBGWBFULL_delay;
wire C405DCRREAD_delay;
wire C405DCRWRITE_delay;
wire C405JTGCAPTUREDR_delay;
wire C405JTGEXTEST_delay;
wire C405JTGPGMOUT_delay;
wire C405JTGSHIFTDR_delay;
wire C405JTGTDO_delay;
wire C405JTGTDOEN_delay;
wire C405JTGUPDATEDR_delay;
wire C405PLBDCUABORT_delay;
wire C405PLBDCUCACHEABLE_delay;
wire C405PLBDCUGUARDED_delay;
wire C405PLBDCUREQUEST_delay;
wire C405PLBDCURNW_delay;
wire C405PLBDCUSIZE2_delay;
wire C405PLBDCUU0ATTR_delay;
wire C405PLBDCUWRITETHRU_delay;
wire C405PLBICUABORT_delay;
wire C405PLBICUCACHEABLE_delay;
wire C405PLBICUREQUEST_delay;
wire C405PLBICUU0ATTR_delay;
wire C405RSTCHIPRESETREQ_delay;
wire C405RSTCORERESETREQ_delay;
wire C405RSTSYSRESETREQ_delay;
wire C405TRCCYCLE_delay;
wire C405TRCTRIGGEREVENTOUT_delay;
wire C405XXXMACHINECHECK_delay;
wire DSOCMBRAMEN_delay;
wire DSOCMBUSY_delay;
wire ISOCMBRAMEN_delay;
wire ISOCMBRAMEVENWRITEEN_delay;
wire ISOCMBRAMODDWRITEEN_delay;

buf (C405CPMCORESLEEPREQ, C405CPMCORESLEEPREQ_delay);
buf (C405CPMMSRCE, C405CPMMSRCE_delay);
buf (C405CPMMSREE, C405CPMMSREE_delay);
buf (C405CPMTIMERIRQ, C405CPMTIMERIRQ_delay);
buf (C405CPMTIMERRESETREQ, C405CPMTIMERRESETREQ_delay);
buf (C405DBGMSRWE, C405DBGMSRWE_delay);
buf (C405DBGSTOPACK, C405DBGSTOPACK_delay);
buf (C405DBGWBCOMPLETE, C405DBGWBCOMPLETE_delay);
buf (C405DBGWBFULL, C405DBGWBFULL_delay);
buf (C405DBGWBIAR[0], C405DBGWBIAR_delay[0]);
buf (C405DBGWBIAR[1], C405DBGWBIAR_delay[1]);
buf (C405DBGWBIAR[2], C405DBGWBIAR_delay[2]);
buf (C405DBGWBIAR[3], C405DBGWBIAR_delay[3]);
buf (C405DBGWBIAR[4], C405DBGWBIAR_delay[4]);
buf (C405DBGWBIAR[5], C405DBGWBIAR_delay[5]);
buf (C405DBGWBIAR[6], C405DBGWBIAR_delay[6]);
buf (C405DBGWBIAR[7], C405DBGWBIAR_delay[7]);
buf (C405DBGWBIAR[8], C405DBGWBIAR_delay[8]);
buf (C405DBGWBIAR[9], C405DBGWBIAR_delay[9]);
buf (C405DBGWBIAR[10], C405DBGWBIAR_delay[10]);
buf (C405DBGWBIAR[11], C405DBGWBIAR_delay[11]);
buf (C405DBGWBIAR[12], C405DBGWBIAR_delay[12]);
buf (C405DBGWBIAR[13], C405DBGWBIAR_delay[13]);
buf (C405DBGWBIAR[14], C405DBGWBIAR_delay[14]);
buf (C405DBGWBIAR[15], C405DBGWBIAR_delay[15]);
buf (C405DBGWBIAR[16], C405DBGWBIAR_delay[16]);
buf (C405DBGWBIAR[17], C405DBGWBIAR_delay[17]);
buf (C405DBGWBIAR[18], C405DBGWBIAR_delay[18]);
buf (C405DBGWBIAR[19], C405DBGWBIAR_delay[19]);
buf (C405DBGWBIAR[20], C405DBGWBIAR_delay[20]);
buf (C405DBGWBIAR[21], C405DBGWBIAR_delay[21]);
buf (C405DBGWBIAR[22], C405DBGWBIAR_delay[22]);
buf (C405DBGWBIAR[23], C405DBGWBIAR_delay[23]);
buf (C405DBGWBIAR[24], C405DBGWBIAR_delay[24]);
buf (C405DBGWBIAR[25], C405DBGWBIAR_delay[25]);
buf (C405DBGWBIAR[26], C405DBGWBIAR_delay[26]);
buf (C405DBGWBIAR[27], C405DBGWBIAR_delay[27]);
buf (C405DBGWBIAR[28], C405DBGWBIAR_delay[28]);
buf (C405DBGWBIAR[29], C405DBGWBIAR_delay[29]);
buf (C405DCRABUS[0], C405DCRABUS_delay[0]);
buf (C405DCRABUS[1], C405DCRABUS_delay[1]);
buf (C405DCRABUS[2], C405DCRABUS_delay[2]);
buf (C405DCRABUS[3], C405DCRABUS_delay[3]);
buf (C405DCRABUS[4], C405DCRABUS_delay[4]);
buf (C405DCRABUS[5], C405DCRABUS_delay[5]);
buf (C405DCRABUS[6], C405DCRABUS_delay[6]);
buf (C405DCRABUS[7], C405DCRABUS_delay[7]);
buf (C405DCRABUS[8], C405DCRABUS_delay[8]);
buf (C405DCRABUS[9], C405DCRABUS_delay[9]);
buf (C405DCRDBUSOUT[0], C405DCRDBUSOUT_delay[0]);
buf (C405DCRDBUSOUT[1], C405DCRDBUSOUT_delay[1]);
buf (C405DCRDBUSOUT[2], C405DCRDBUSOUT_delay[2]);
buf (C405DCRDBUSOUT[3], C405DCRDBUSOUT_delay[3]);
buf (C405DCRDBUSOUT[4], C405DCRDBUSOUT_delay[4]);
buf (C405DCRDBUSOUT[5], C405DCRDBUSOUT_delay[5]);
buf (C405DCRDBUSOUT[6], C405DCRDBUSOUT_delay[6]);
buf (C405DCRDBUSOUT[7], C405DCRDBUSOUT_delay[7]);
buf (C405DCRDBUSOUT[8], C405DCRDBUSOUT_delay[8]);
buf (C405DCRDBUSOUT[9], C405DCRDBUSOUT_delay[9]);
buf (C405DCRDBUSOUT[10], C405DCRDBUSOUT_delay[10]);
buf (C405DCRDBUSOUT[11], C405DCRDBUSOUT_delay[11]);
buf (C405DCRDBUSOUT[12], C405DCRDBUSOUT_delay[12]);
buf (C405DCRDBUSOUT[13], C405DCRDBUSOUT_delay[13]);
buf (C405DCRDBUSOUT[14], C405DCRDBUSOUT_delay[14]);
buf (C405DCRDBUSOUT[15], C405DCRDBUSOUT_delay[15]);
buf (C405DCRDBUSOUT[16], C405DCRDBUSOUT_delay[16]);
buf (C405DCRDBUSOUT[17], C405DCRDBUSOUT_delay[17]);
buf (C405DCRDBUSOUT[18], C405DCRDBUSOUT_delay[18]);
buf (C405DCRDBUSOUT[19], C405DCRDBUSOUT_delay[19]);
buf (C405DCRDBUSOUT[20], C405DCRDBUSOUT_delay[20]);
buf (C405DCRDBUSOUT[21], C405DCRDBUSOUT_delay[21]);
buf (C405DCRDBUSOUT[22], C405DCRDBUSOUT_delay[22]);
buf (C405DCRDBUSOUT[23], C405DCRDBUSOUT_delay[23]);
buf (C405DCRDBUSOUT[24], C405DCRDBUSOUT_delay[24]);
buf (C405DCRDBUSOUT[25], C405DCRDBUSOUT_delay[25]);
buf (C405DCRDBUSOUT[26], C405DCRDBUSOUT_delay[26]);
buf (C405DCRDBUSOUT[27], C405DCRDBUSOUT_delay[27]);
buf (C405DCRDBUSOUT[28], C405DCRDBUSOUT_delay[28]);
buf (C405DCRDBUSOUT[29], C405DCRDBUSOUT_delay[29]);
buf (C405DCRDBUSOUT[30], C405DCRDBUSOUT_delay[30]);
buf (C405DCRDBUSOUT[31], C405DCRDBUSOUT_delay[31]);
buf (C405DCRREAD, C405DCRREAD_delay);
buf (C405DCRWRITE, C405DCRWRITE_delay);
buf (C405JTGCAPTUREDR, C405JTGCAPTUREDR_delay);
buf (C405JTGEXTEST, C405JTGEXTEST_delay);
buf (C405JTGPGMOUT, C405JTGPGMOUT_delay);
buf (C405JTGSHIFTDR, C405JTGSHIFTDR_delay);
buf (C405JTGTDO, C405JTGTDO_delay);
buf (C405JTGTDOEN, C405JTGTDOEN_delay);
buf (C405JTGUPDATEDR, C405JTGUPDATEDR_delay);
buf (C405PLBDCUABORT, C405PLBDCUABORT_delay);
buf (C405PLBDCUABUS[0], C405PLBDCUABUS_delay[0]);
buf (C405PLBDCUABUS[1], C405PLBDCUABUS_delay[1]);
buf (C405PLBDCUABUS[2], C405PLBDCUABUS_delay[2]);
buf (C405PLBDCUABUS[3], C405PLBDCUABUS_delay[3]);
buf (C405PLBDCUABUS[4], C405PLBDCUABUS_delay[4]);
buf (C405PLBDCUABUS[5], C405PLBDCUABUS_delay[5]);
buf (C405PLBDCUABUS[6], C405PLBDCUABUS_delay[6]);
buf (C405PLBDCUABUS[7], C405PLBDCUABUS_delay[7]);
buf (C405PLBDCUABUS[8], C405PLBDCUABUS_delay[8]);
buf (C405PLBDCUABUS[9], C405PLBDCUABUS_delay[9]);
buf (C405PLBDCUABUS[10], C405PLBDCUABUS_delay[10]);
buf (C405PLBDCUABUS[11], C405PLBDCUABUS_delay[11]);
buf (C405PLBDCUABUS[12], C405PLBDCUABUS_delay[12]);
buf (C405PLBDCUABUS[13], C405PLBDCUABUS_delay[13]);
buf (C405PLBDCUABUS[14], C405PLBDCUABUS_delay[14]);
buf (C405PLBDCUABUS[15], C405PLBDCUABUS_delay[15]);
buf (C405PLBDCUABUS[16], C405PLBDCUABUS_delay[16]);
buf (C405PLBDCUABUS[17], C405PLBDCUABUS_delay[17]);
buf (C405PLBDCUABUS[18], C405PLBDCUABUS_delay[18]);
buf (C405PLBDCUABUS[19], C405PLBDCUABUS_delay[19]);
buf (C405PLBDCUABUS[20], C405PLBDCUABUS_delay[20]);
buf (C405PLBDCUABUS[21], C405PLBDCUABUS_delay[21]);
buf (C405PLBDCUABUS[22], C405PLBDCUABUS_delay[22]);
buf (C405PLBDCUABUS[23], C405PLBDCUABUS_delay[23]);
buf (C405PLBDCUABUS[24], C405PLBDCUABUS_delay[24]);
buf (C405PLBDCUABUS[25], C405PLBDCUABUS_delay[25]);
buf (C405PLBDCUABUS[26], C405PLBDCUABUS_delay[26]);
buf (C405PLBDCUABUS[27], C405PLBDCUABUS_delay[27]);
buf (C405PLBDCUABUS[28], C405PLBDCUABUS_delay[28]);
buf (C405PLBDCUABUS[29], C405PLBDCUABUS_delay[29]);
buf (C405PLBDCUABUS[30], C405PLBDCUABUS_delay[30]);
buf (C405PLBDCUABUS[31], C405PLBDCUABUS_delay[31]);
buf (C405PLBDCUBE[0], C405PLBDCUBE_delay[0]);
buf (C405PLBDCUBE[1], C405PLBDCUBE_delay[1]);
buf (C405PLBDCUBE[2], C405PLBDCUBE_delay[2]);
buf (C405PLBDCUBE[3], C405PLBDCUBE_delay[3]);
buf (C405PLBDCUBE[4], C405PLBDCUBE_delay[4]);
buf (C405PLBDCUBE[5], C405PLBDCUBE_delay[5]);
buf (C405PLBDCUBE[6], C405PLBDCUBE_delay[6]);
buf (C405PLBDCUBE[7], C405PLBDCUBE_delay[7]);
buf (C405PLBDCUCACHEABLE, C405PLBDCUCACHEABLE_delay);
buf (C405PLBDCUGUARDED, C405PLBDCUGUARDED_delay);
buf (C405PLBDCUPRIORITY[0], C405PLBDCUPRIORITY_delay[0]);
buf (C405PLBDCUPRIORITY[1], C405PLBDCUPRIORITY_delay[1]);
buf (C405PLBDCUREQUEST, C405PLBDCUREQUEST_delay);
buf (C405PLBDCURNW, C405PLBDCURNW_delay);
buf (C405PLBDCUSIZE2, C405PLBDCUSIZE2_delay);
buf (C405PLBDCUU0ATTR, C405PLBDCUU0ATTR_delay);
buf (C405PLBDCUWRDBUS[0], C405PLBDCUWRDBUS_delay[0]);
buf (C405PLBDCUWRDBUS[1], C405PLBDCUWRDBUS_delay[1]);
buf (C405PLBDCUWRDBUS[2], C405PLBDCUWRDBUS_delay[2]);
buf (C405PLBDCUWRDBUS[3], C405PLBDCUWRDBUS_delay[3]);
buf (C405PLBDCUWRDBUS[4], C405PLBDCUWRDBUS_delay[4]);
buf (C405PLBDCUWRDBUS[5], C405PLBDCUWRDBUS_delay[5]);
buf (C405PLBDCUWRDBUS[6], C405PLBDCUWRDBUS_delay[6]);
buf (C405PLBDCUWRDBUS[7], C405PLBDCUWRDBUS_delay[7]);
buf (C405PLBDCUWRDBUS[8], C405PLBDCUWRDBUS_delay[8]);
buf (C405PLBDCUWRDBUS[9], C405PLBDCUWRDBUS_delay[9]);
buf (C405PLBDCUWRDBUS[10], C405PLBDCUWRDBUS_delay[10]);
buf (C405PLBDCUWRDBUS[11], C405PLBDCUWRDBUS_delay[11]);
buf (C405PLBDCUWRDBUS[12], C405PLBDCUWRDBUS_delay[12]);
buf (C405PLBDCUWRDBUS[13], C405PLBDCUWRDBUS_delay[13]);
buf (C405PLBDCUWRDBUS[14], C405PLBDCUWRDBUS_delay[14]);
buf (C405PLBDCUWRDBUS[15], C405PLBDCUWRDBUS_delay[15]);
buf (C405PLBDCUWRDBUS[16], C405PLBDCUWRDBUS_delay[16]);
buf (C405PLBDCUWRDBUS[17], C405PLBDCUWRDBUS_delay[17]);
buf (C405PLBDCUWRDBUS[18], C405PLBDCUWRDBUS_delay[18]);
buf (C405PLBDCUWRDBUS[19], C405PLBDCUWRDBUS_delay[19]);
buf (C405PLBDCUWRDBUS[20], C405PLBDCUWRDBUS_delay[20]);
buf (C405PLBDCUWRDBUS[21], C405PLBDCUWRDBUS_delay[21]);
buf (C405PLBDCUWRDBUS[22], C405PLBDCUWRDBUS_delay[22]);
buf (C405PLBDCUWRDBUS[23], C405PLBDCUWRDBUS_delay[23]);
buf (C405PLBDCUWRDBUS[24], C405PLBDCUWRDBUS_delay[24]);
buf (C405PLBDCUWRDBUS[25], C405PLBDCUWRDBUS_delay[25]);
buf (C405PLBDCUWRDBUS[26], C405PLBDCUWRDBUS_delay[26]);
buf (C405PLBDCUWRDBUS[27], C405PLBDCUWRDBUS_delay[27]);
buf (C405PLBDCUWRDBUS[28], C405PLBDCUWRDBUS_delay[28]);
buf (C405PLBDCUWRDBUS[29], C405PLBDCUWRDBUS_delay[29]);
buf (C405PLBDCUWRDBUS[30], C405PLBDCUWRDBUS_delay[30]);
buf (C405PLBDCUWRDBUS[31], C405PLBDCUWRDBUS_delay[31]);
buf (C405PLBDCUWRDBUS[32], C405PLBDCUWRDBUS_delay[32]);
buf (C405PLBDCUWRDBUS[33], C405PLBDCUWRDBUS_delay[33]);
buf (C405PLBDCUWRDBUS[34], C405PLBDCUWRDBUS_delay[34]);
buf (C405PLBDCUWRDBUS[35], C405PLBDCUWRDBUS_delay[35]);
buf (C405PLBDCUWRDBUS[36], C405PLBDCUWRDBUS_delay[36]);
buf (C405PLBDCUWRDBUS[37], C405PLBDCUWRDBUS_delay[37]);
buf (C405PLBDCUWRDBUS[38], C405PLBDCUWRDBUS_delay[38]);
buf (C405PLBDCUWRDBUS[39], C405PLBDCUWRDBUS_delay[39]);
buf (C405PLBDCUWRDBUS[40], C405PLBDCUWRDBUS_delay[40]);
buf (C405PLBDCUWRDBUS[41], C405PLBDCUWRDBUS_delay[41]);
buf (C405PLBDCUWRDBUS[42], C405PLBDCUWRDBUS_delay[42]);
buf (C405PLBDCUWRDBUS[43], C405PLBDCUWRDBUS_delay[43]);
buf (C405PLBDCUWRDBUS[44], C405PLBDCUWRDBUS_delay[44]);
buf (C405PLBDCUWRDBUS[45], C405PLBDCUWRDBUS_delay[45]);
buf (C405PLBDCUWRDBUS[46], C405PLBDCUWRDBUS_delay[46]);
buf (C405PLBDCUWRDBUS[47], C405PLBDCUWRDBUS_delay[47]);
buf (C405PLBDCUWRDBUS[48], C405PLBDCUWRDBUS_delay[48]);
buf (C405PLBDCUWRDBUS[49], C405PLBDCUWRDBUS_delay[49]);
buf (C405PLBDCUWRDBUS[50], C405PLBDCUWRDBUS_delay[50]);
buf (C405PLBDCUWRDBUS[51], C405PLBDCUWRDBUS_delay[51]);
buf (C405PLBDCUWRDBUS[52], C405PLBDCUWRDBUS_delay[52]);
buf (C405PLBDCUWRDBUS[53], C405PLBDCUWRDBUS_delay[53]);
buf (C405PLBDCUWRDBUS[54], C405PLBDCUWRDBUS_delay[54]);
buf (C405PLBDCUWRDBUS[55], C405PLBDCUWRDBUS_delay[55]);
buf (C405PLBDCUWRDBUS[56], C405PLBDCUWRDBUS_delay[56]);
buf (C405PLBDCUWRDBUS[57], C405PLBDCUWRDBUS_delay[57]);
buf (C405PLBDCUWRDBUS[58], C405PLBDCUWRDBUS_delay[58]);
buf (C405PLBDCUWRDBUS[59], C405PLBDCUWRDBUS_delay[59]);
buf (C405PLBDCUWRDBUS[60], C405PLBDCUWRDBUS_delay[60]);
buf (C405PLBDCUWRDBUS[61], C405PLBDCUWRDBUS_delay[61]);
buf (C405PLBDCUWRDBUS[62], C405PLBDCUWRDBUS_delay[62]);
buf (C405PLBDCUWRDBUS[63], C405PLBDCUWRDBUS_delay[63]);
buf (C405PLBDCUWRITETHRU, C405PLBDCUWRITETHRU_delay);
buf (C405PLBICUABORT, C405PLBICUABORT_delay);
buf (C405PLBICUABUS[0], C405PLBICUABUS_delay[0]);
buf (C405PLBICUABUS[1], C405PLBICUABUS_delay[1]);
buf (C405PLBICUABUS[2], C405PLBICUABUS_delay[2]);
buf (C405PLBICUABUS[3], C405PLBICUABUS_delay[3]);
buf (C405PLBICUABUS[4], C405PLBICUABUS_delay[4]);
buf (C405PLBICUABUS[5], C405PLBICUABUS_delay[5]);
buf (C405PLBICUABUS[6], C405PLBICUABUS_delay[6]);
buf (C405PLBICUABUS[7], C405PLBICUABUS_delay[7]);
buf (C405PLBICUABUS[8], C405PLBICUABUS_delay[8]);
buf (C405PLBICUABUS[9], C405PLBICUABUS_delay[9]);
buf (C405PLBICUABUS[10], C405PLBICUABUS_delay[10]);
buf (C405PLBICUABUS[11], C405PLBICUABUS_delay[11]);
buf (C405PLBICUABUS[12], C405PLBICUABUS_delay[12]);
buf (C405PLBICUABUS[13], C405PLBICUABUS_delay[13]);
buf (C405PLBICUABUS[14], C405PLBICUABUS_delay[14]);
buf (C405PLBICUABUS[15], C405PLBICUABUS_delay[15]);
buf (C405PLBICUABUS[16], C405PLBICUABUS_delay[16]);
buf (C405PLBICUABUS[17], C405PLBICUABUS_delay[17]);
buf (C405PLBICUABUS[18], C405PLBICUABUS_delay[18]);
buf (C405PLBICUABUS[19], C405PLBICUABUS_delay[19]);
buf (C405PLBICUABUS[20], C405PLBICUABUS_delay[20]);
buf (C405PLBICUABUS[21], C405PLBICUABUS_delay[21]);
buf (C405PLBICUABUS[22], C405PLBICUABUS_delay[22]);
buf (C405PLBICUABUS[23], C405PLBICUABUS_delay[23]);
buf (C405PLBICUABUS[24], C405PLBICUABUS_delay[24]);
buf (C405PLBICUABUS[25], C405PLBICUABUS_delay[25]);
buf (C405PLBICUABUS[26], C405PLBICUABUS_delay[26]);
buf (C405PLBICUABUS[27], C405PLBICUABUS_delay[27]);
buf (C405PLBICUABUS[28], C405PLBICUABUS_delay[28]);
buf (C405PLBICUABUS[29], C405PLBICUABUS_delay[29]);
buf (C405PLBICUCACHEABLE, C405PLBICUCACHEABLE_delay);
buf (C405PLBICUPRIORITY[0], C405PLBICUPRIORITY_delay[0]);
buf (C405PLBICUPRIORITY[1], C405PLBICUPRIORITY_delay[1]);
buf (C405PLBICUREQUEST, C405PLBICUREQUEST_delay);
buf (C405PLBICUSIZE[2], C405PLBICUSIZE_delay[2]);
buf (C405PLBICUSIZE[3], C405PLBICUSIZE_delay[3]);
buf (C405PLBICUU0ATTR, C405PLBICUU0ATTR_delay);
buf (C405RSTCHIPRESETREQ, C405RSTCHIPRESETREQ_delay);
buf (C405RSTCORERESETREQ, C405RSTCORERESETREQ_delay);
buf (C405RSTSYSRESETREQ, C405RSTSYSRESETREQ_delay);
buf (C405TRCCYCLE, C405TRCCYCLE_delay);
buf (C405TRCEVENEXECUTIONSTATUS[0], C405TRCEVENEXECUTIONSTATUS_delay[0]);
buf (C405TRCEVENEXECUTIONSTATUS[1], C405TRCEVENEXECUTIONSTATUS_delay[1]);
buf (C405TRCODDEXECUTIONSTATUS[0], C405TRCODDEXECUTIONSTATUS_delay[0]);
buf (C405TRCODDEXECUTIONSTATUS[1], C405TRCODDEXECUTIONSTATUS_delay[1]);
buf (C405TRCTRACESTATUS[0], C405TRCTRACESTATUS_delay[0]);
buf (C405TRCTRACESTATUS[1], C405TRCTRACESTATUS_delay[1]);
buf (C405TRCTRACESTATUS[2], C405TRCTRACESTATUS_delay[2]);
buf (C405TRCTRACESTATUS[3], C405TRCTRACESTATUS_delay[3]);
buf (C405TRCTRIGGEREVENTOUT, C405TRCTRIGGEREVENTOUT_delay);
buf (C405TRCTRIGGEREVENTTYPE[0], C405TRCTRIGGEREVENTTYPE_delay[0]);
buf (C405TRCTRIGGEREVENTTYPE[1], C405TRCTRIGGEREVENTTYPE_delay[1]);
buf (C405TRCTRIGGEREVENTTYPE[2], C405TRCTRIGGEREVENTTYPE_delay[2]);
buf (C405TRCTRIGGEREVENTTYPE[3], C405TRCTRIGGEREVENTTYPE_delay[3]);
buf (C405TRCTRIGGEREVENTTYPE[4], C405TRCTRIGGEREVENTTYPE_delay[4]);
buf (C405TRCTRIGGEREVENTTYPE[5], C405TRCTRIGGEREVENTTYPE_delay[5]);
buf (C405TRCTRIGGEREVENTTYPE[6], C405TRCTRIGGEREVENTTYPE_delay[6]);
buf (C405TRCTRIGGEREVENTTYPE[7], C405TRCTRIGGEREVENTTYPE_delay[7]);
buf (C405TRCTRIGGEREVENTTYPE[8], C405TRCTRIGGEREVENTTYPE_delay[8]);
buf (C405TRCTRIGGEREVENTTYPE[9], C405TRCTRIGGEREVENTTYPE_delay[9]);
buf (C405TRCTRIGGEREVENTTYPE[10], C405TRCTRIGGEREVENTTYPE_delay[10]);
buf (C405XXXMACHINECHECK, C405XXXMACHINECHECK_delay);
buf (DSOCMBRAMABUS[8], DSOCMBRAMABUS_delay[8]);
buf (DSOCMBRAMABUS[9], DSOCMBRAMABUS_delay[9]);
buf (DSOCMBRAMABUS[10], DSOCMBRAMABUS_delay[10]);
buf (DSOCMBRAMABUS[11], DSOCMBRAMABUS_delay[11]);
buf (DSOCMBRAMABUS[12], DSOCMBRAMABUS_delay[12]);
buf (DSOCMBRAMABUS[13], DSOCMBRAMABUS_delay[13]);
buf (DSOCMBRAMABUS[14], DSOCMBRAMABUS_delay[14]);
buf (DSOCMBRAMABUS[15], DSOCMBRAMABUS_delay[15]);
buf (DSOCMBRAMABUS[16], DSOCMBRAMABUS_delay[16]);
buf (DSOCMBRAMABUS[17], DSOCMBRAMABUS_delay[17]);
buf (DSOCMBRAMABUS[18], DSOCMBRAMABUS_delay[18]);
buf (DSOCMBRAMABUS[19], DSOCMBRAMABUS_delay[19]);
buf (DSOCMBRAMABUS[20], DSOCMBRAMABUS_delay[20]);
buf (DSOCMBRAMABUS[21], DSOCMBRAMABUS_delay[21]);
buf (DSOCMBRAMABUS[22], DSOCMBRAMABUS_delay[22]);
buf (DSOCMBRAMABUS[23], DSOCMBRAMABUS_delay[23]);
buf (DSOCMBRAMABUS[24], DSOCMBRAMABUS_delay[24]);
buf (DSOCMBRAMABUS[25], DSOCMBRAMABUS_delay[25]);
buf (DSOCMBRAMABUS[26], DSOCMBRAMABUS_delay[26]);
buf (DSOCMBRAMABUS[27], DSOCMBRAMABUS_delay[27]);
buf (DSOCMBRAMABUS[28], DSOCMBRAMABUS_delay[28]);
buf (DSOCMBRAMABUS[29], DSOCMBRAMABUS_delay[29]);
buf (DSOCMBRAMBYTEWRITE[0], DSOCMBRAMBYTEWRITE_delay[0]);
buf (DSOCMBRAMBYTEWRITE[1], DSOCMBRAMBYTEWRITE_delay[1]);
buf (DSOCMBRAMBYTEWRITE[2], DSOCMBRAMBYTEWRITE_delay[2]);
buf (DSOCMBRAMBYTEWRITE[3], DSOCMBRAMBYTEWRITE_delay[3]);
buf (DSOCMBRAMEN, DSOCMBRAMEN_delay);
buf (DSOCMBRAMWRDBUS[0], DSOCMBRAMWRDBUS_delay[0]);
buf (DSOCMBRAMWRDBUS[1], DSOCMBRAMWRDBUS_delay[1]);
buf (DSOCMBRAMWRDBUS[2], DSOCMBRAMWRDBUS_delay[2]);
buf (DSOCMBRAMWRDBUS[3], DSOCMBRAMWRDBUS_delay[3]);
buf (DSOCMBRAMWRDBUS[4], DSOCMBRAMWRDBUS_delay[4]);
buf (DSOCMBRAMWRDBUS[5], DSOCMBRAMWRDBUS_delay[5]);
buf (DSOCMBRAMWRDBUS[6], DSOCMBRAMWRDBUS_delay[6]);
buf (DSOCMBRAMWRDBUS[7], DSOCMBRAMWRDBUS_delay[7]);
buf (DSOCMBRAMWRDBUS[8], DSOCMBRAMWRDBUS_delay[8]);
buf (DSOCMBRAMWRDBUS[9], DSOCMBRAMWRDBUS_delay[9]);
buf (DSOCMBRAMWRDBUS[10], DSOCMBRAMWRDBUS_delay[10]);
buf (DSOCMBRAMWRDBUS[11], DSOCMBRAMWRDBUS_delay[11]);
buf (DSOCMBRAMWRDBUS[12], DSOCMBRAMWRDBUS_delay[12]);
buf (DSOCMBRAMWRDBUS[13], DSOCMBRAMWRDBUS_delay[13]);
buf (DSOCMBRAMWRDBUS[14], DSOCMBRAMWRDBUS_delay[14]);
buf (DSOCMBRAMWRDBUS[15], DSOCMBRAMWRDBUS_delay[15]);
buf (DSOCMBRAMWRDBUS[16], DSOCMBRAMWRDBUS_delay[16]);
buf (DSOCMBRAMWRDBUS[17], DSOCMBRAMWRDBUS_delay[17]);
buf (DSOCMBRAMWRDBUS[18], DSOCMBRAMWRDBUS_delay[18]);
buf (DSOCMBRAMWRDBUS[19], DSOCMBRAMWRDBUS_delay[19]);
buf (DSOCMBRAMWRDBUS[20], DSOCMBRAMWRDBUS_delay[20]);
buf (DSOCMBRAMWRDBUS[21], DSOCMBRAMWRDBUS_delay[21]);
buf (DSOCMBRAMWRDBUS[22], DSOCMBRAMWRDBUS_delay[22]);
buf (DSOCMBRAMWRDBUS[23], DSOCMBRAMWRDBUS_delay[23]);
buf (DSOCMBRAMWRDBUS[24], DSOCMBRAMWRDBUS_delay[24]);
buf (DSOCMBRAMWRDBUS[25], DSOCMBRAMWRDBUS_delay[25]);
buf (DSOCMBRAMWRDBUS[26], DSOCMBRAMWRDBUS_delay[26]);
buf (DSOCMBRAMWRDBUS[27], DSOCMBRAMWRDBUS_delay[27]);
buf (DSOCMBRAMWRDBUS[28], DSOCMBRAMWRDBUS_delay[28]);
buf (DSOCMBRAMWRDBUS[29], DSOCMBRAMWRDBUS_delay[29]);
buf (DSOCMBRAMWRDBUS[30], DSOCMBRAMWRDBUS_delay[30]);
buf (DSOCMBRAMWRDBUS[31], DSOCMBRAMWRDBUS_delay[31]);
buf (DSOCMBUSY, DSOCMBUSY_delay);
buf (ISOCMBRAMEN, ISOCMBRAMEN_delay);
buf (ISOCMBRAMEVENWRITEEN, ISOCMBRAMEVENWRITEEN_delay);
buf (ISOCMBRAMODDWRITEEN, ISOCMBRAMODDWRITEEN_delay);
buf (ISOCMBRAMRDABUS[8], ISOCMBRAMRDABUS_delay[8]);
buf (ISOCMBRAMRDABUS[9], ISOCMBRAMRDABUS_delay[9]);
buf (ISOCMBRAMRDABUS[10], ISOCMBRAMRDABUS_delay[10]);
buf (ISOCMBRAMRDABUS[11], ISOCMBRAMRDABUS_delay[11]);
buf (ISOCMBRAMRDABUS[12], ISOCMBRAMRDABUS_delay[12]);
buf (ISOCMBRAMRDABUS[13], ISOCMBRAMRDABUS_delay[13]);
buf (ISOCMBRAMRDABUS[14], ISOCMBRAMRDABUS_delay[14]);
buf (ISOCMBRAMRDABUS[15], ISOCMBRAMRDABUS_delay[15]);
buf (ISOCMBRAMRDABUS[16], ISOCMBRAMRDABUS_delay[16]);
buf (ISOCMBRAMRDABUS[17], ISOCMBRAMRDABUS_delay[17]);
buf (ISOCMBRAMRDABUS[18], ISOCMBRAMRDABUS_delay[18]);
buf (ISOCMBRAMRDABUS[19], ISOCMBRAMRDABUS_delay[19]);
buf (ISOCMBRAMRDABUS[20], ISOCMBRAMRDABUS_delay[20]);
buf (ISOCMBRAMRDABUS[21], ISOCMBRAMRDABUS_delay[21]);
buf (ISOCMBRAMRDABUS[22], ISOCMBRAMRDABUS_delay[22]);
buf (ISOCMBRAMRDABUS[23], ISOCMBRAMRDABUS_delay[23]);
buf (ISOCMBRAMRDABUS[24], ISOCMBRAMRDABUS_delay[24]);
buf (ISOCMBRAMRDABUS[25], ISOCMBRAMRDABUS_delay[25]);
buf (ISOCMBRAMRDABUS[26], ISOCMBRAMRDABUS_delay[26]);
buf (ISOCMBRAMRDABUS[27], ISOCMBRAMRDABUS_delay[27]);
buf (ISOCMBRAMRDABUS[28], ISOCMBRAMRDABUS_delay[28]);
buf (ISOCMBRAMWRABUS[8], ISOCMBRAMWRABUS_delay[8]);
buf (ISOCMBRAMWRABUS[9], ISOCMBRAMWRABUS_delay[9]);
buf (ISOCMBRAMWRABUS[10], ISOCMBRAMWRABUS_delay[10]);
buf (ISOCMBRAMWRABUS[11], ISOCMBRAMWRABUS_delay[11]);
buf (ISOCMBRAMWRABUS[12], ISOCMBRAMWRABUS_delay[12]);
buf (ISOCMBRAMWRABUS[13], ISOCMBRAMWRABUS_delay[13]);
buf (ISOCMBRAMWRABUS[14], ISOCMBRAMWRABUS_delay[14]);
buf (ISOCMBRAMWRABUS[15], ISOCMBRAMWRABUS_delay[15]);
buf (ISOCMBRAMWRABUS[16], ISOCMBRAMWRABUS_delay[16]);
buf (ISOCMBRAMWRABUS[17], ISOCMBRAMWRABUS_delay[17]);
buf (ISOCMBRAMWRABUS[18], ISOCMBRAMWRABUS_delay[18]);
buf (ISOCMBRAMWRABUS[19], ISOCMBRAMWRABUS_delay[19]);
buf (ISOCMBRAMWRABUS[20], ISOCMBRAMWRABUS_delay[20]);
buf (ISOCMBRAMWRABUS[21], ISOCMBRAMWRABUS_delay[21]);
buf (ISOCMBRAMWRABUS[22], ISOCMBRAMWRABUS_delay[22]);
buf (ISOCMBRAMWRABUS[23], ISOCMBRAMWRABUS_delay[23]);
buf (ISOCMBRAMWRABUS[24], ISOCMBRAMWRABUS_delay[24]);
buf (ISOCMBRAMWRABUS[25], ISOCMBRAMWRABUS_delay[25]);
buf (ISOCMBRAMWRABUS[26], ISOCMBRAMWRABUS_delay[26]);
buf (ISOCMBRAMWRABUS[27], ISOCMBRAMWRABUS_delay[27]);
buf (ISOCMBRAMWRABUS[28], ISOCMBRAMWRABUS_delay[28]);
buf (ISOCMBRAMWRDBUS[0], ISOCMBRAMWRDBUS_delay[0]);
buf (ISOCMBRAMWRDBUS[1], ISOCMBRAMWRDBUS_delay[1]);
buf (ISOCMBRAMWRDBUS[2], ISOCMBRAMWRDBUS_delay[2]);
buf (ISOCMBRAMWRDBUS[3], ISOCMBRAMWRDBUS_delay[3]);
buf (ISOCMBRAMWRDBUS[4], ISOCMBRAMWRDBUS_delay[4]);
buf (ISOCMBRAMWRDBUS[5], ISOCMBRAMWRDBUS_delay[5]);
buf (ISOCMBRAMWRDBUS[6], ISOCMBRAMWRDBUS_delay[6]);
buf (ISOCMBRAMWRDBUS[7], ISOCMBRAMWRDBUS_delay[7]);
buf (ISOCMBRAMWRDBUS[8], ISOCMBRAMWRDBUS_delay[8]);
buf (ISOCMBRAMWRDBUS[9], ISOCMBRAMWRDBUS_delay[9]);
buf (ISOCMBRAMWRDBUS[10], ISOCMBRAMWRDBUS_delay[10]);
buf (ISOCMBRAMWRDBUS[11], ISOCMBRAMWRDBUS_delay[11]);
buf (ISOCMBRAMWRDBUS[12], ISOCMBRAMWRDBUS_delay[12]);
buf (ISOCMBRAMWRDBUS[13], ISOCMBRAMWRDBUS_delay[13]);
buf (ISOCMBRAMWRDBUS[14], ISOCMBRAMWRDBUS_delay[14]);
buf (ISOCMBRAMWRDBUS[15], ISOCMBRAMWRDBUS_delay[15]);
buf (ISOCMBRAMWRDBUS[16], ISOCMBRAMWRDBUS_delay[16]);
buf (ISOCMBRAMWRDBUS[17], ISOCMBRAMWRDBUS_delay[17]);
buf (ISOCMBRAMWRDBUS[18], ISOCMBRAMWRDBUS_delay[18]);
buf (ISOCMBRAMWRDBUS[19], ISOCMBRAMWRDBUS_delay[19]);
buf (ISOCMBRAMWRDBUS[20], ISOCMBRAMWRDBUS_delay[20]);
buf (ISOCMBRAMWRDBUS[21], ISOCMBRAMWRDBUS_delay[21]);
buf (ISOCMBRAMWRDBUS[22], ISOCMBRAMWRDBUS_delay[22]);
buf (ISOCMBRAMWRDBUS[23], ISOCMBRAMWRDBUS_delay[23]);
buf (ISOCMBRAMWRDBUS[24], ISOCMBRAMWRDBUS_delay[24]);
buf (ISOCMBRAMWRDBUS[25], ISOCMBRAMWRDBUS_delay[25]);
buf (ISOCMBRAMWRDBUS[26], ISOCMBRAMWRDBUS_delay[26]);
buf (ISOCMBRAMWRDBUS[27], ISOCMBRAMWRDBUS_delay[27]);
buf (ISOCMBRAMWRDBUS[28], ISOCMBRAMWRDBUS_delay[28]);
buf (ISOCMBRAMWRDBUS[29], ISOCMBRAMWRDBUS_delay[29]);
buf (ISOCMBRAMWRDBUS[30], ISOCMBRAMWRDBUS_delay[30]);
buf (ISOCMBRAMWRDBUS[31], ISOCMBRAMWRDBUS_delay[31]);

buf (BRAMDSOCMCLK_delay, BRAMDSOCMCLK);
buf (BRAMDSOCMRDDBUS_delay[0], BRAMDSOCMRDDBUS[0]);
buf (BRAMDSOCMRDDBUS_delay[1], BRAMDSOCMRDDBUS[1]);
buf (BRAMDSOCMRDDBUS_delay[2], BRAMDSOCMRDDBUS[2]);
buf (BRAMDSOCMRDDBUS_delay[3], BRAMDSOCMRDDBUS[3]);
buf (BRAMDSOCMRDDBUS_delay[4], BRAMDSOCMRDDBUS[4]);
buf (BRAMDSOCMRDDBUS_delay[5], BRAMDSOCMRDDBUS[5]);
buf (BRAMDSOCMRDDBUS_delay[6], BRAMDSOCMRDDBUS[6]);
buf (BRAMDSOCMRDDBUS_delay[7], BRAMDSOCMRDDBUS[7]);
buf (BRAMDSOCMRDDBUS_delay[8], BRAMDSOCMRDDBUS[8]);
buf (BRAMDSOCMRDDBUS_delay[9], BRAMDSOCMRDDBUS[9]);
buf (BRAMDSOCMRDDBUS_delay[10], BRAMDSOCMRDDBUS[10]);
buf (BRAMDSOCMRDDBUS_delay[11], BRAMDSOCMRDDBUS[11]);
buf (BRAMDSOCMRDDBUS_delay[12], BRAMDSOCMRDDBUS[12]);
buf (BRAMDSOCMRDDBUS_delay[13], BRAMDSOCMRDDBUS[13]);
buf (BRAMDSOCMRDDBUS_delay[14], BRAMDSOCMRDDBUS[14]);
buf (BRAMDSOCMRDDBUS_delay[15], BRAMDSOCMRDDBUS[15]);
buf (BRAMDSOCMRDDBUS_delay[16], BRAMDSOCMRDDBUS[16]);
buf (BRAMDSOCMRDDBUS_delay[17], BRAMDSOCMRDDBUS[17]);
buf (BRAMDSOCMRDDBUS_delay[18], BRAMDSOCMRDDBUS[18]);
buf (BRAMDSOCMRDDBUS_delay[19], BRAMDSOCMRDDBUS[19]);
buf (BRAMDSOCMRDDBUS_delay[20], BRAMDSOCMRDDBUS[20]);
buf (BRAMDSOCMRDDBUS_delay[21], BRAMDSOCMRDDBUS[21]);
buf (BRAMDSOCMRDDBUS_delay[22], BRAMDSOCMRDDBUS[22]);
buf (BRAMDSOCMRDDBUS_delay[23], BRAMDSOCMRDDBUS[23]);
buf (BRAMDSOCMRDDBUS_delay[24], BRAMDSOCMRDDBUS[24]);
buf (BRAMDSOCMRDDBUS_delay[25], BRAMDSOCMRDDBUS[25]);
buf (BRAMDSOCMRDDBUS_delay[26], BRAMDSOCMRDDBUS[26]);
buf (BRAMDSOCMRDDBUS_delay[27], BRAMDSOCMRDDBUS[27]);
buf (BRAMDSOCMRDDBUS_delay[28], BRAMDSOCMRDDBUS[28]);
buf (BRAMDSOCMRDDBUS_delay[29], BRAMDSOCMRDDBUS[29]);
buf (BRAMDSOCMRDDBUS_delay[30], BRAMDSOCMRDDBUS[30]);
buf (BRAMDSOCMRDDBUS_delay[31], BRAMDSOCMRDDBUS[31]);
buf (BRAMISOCMCLK_delay, BRAMISOCMCLK);
buf (BRAMISOCMRDDBUS_delay[0], BRAMISOCMRDDBUS[0]);
buf (BRAMISOCMRDDBUS_delay[1], BRAMISOCMRDDBUS[1]);
buf (BRAMISOCMRDDBUS_delay[2], BRAMISOCMRDDBUS[2]);
buf (BRAMISOCMRDDBUS_delay[3], BRAMISOCMRDDBUS[3]);
buf (BRAMISOCMRDDBUS_delay[4], BRAMISOCMRDDBUS[4]);
buf (BRAMISOCMRDDBUS_delay[5], BRAMISOCMRDDBUS[5]);
buf (BRAMISOCMRDDBUS_delay[6], BRAMISOCMRDDBUS[6]);
buf (BRAMISOCMRDDBUS_delay[7], BRAMISOCMRDDBUS[7]);
buf (BRAMISOCMRDDBUS_delay[8], BRAMISOCMRDDBUS[8]);
buf (BRAMISOCMRDDBUS_delay[9], BRAMISOCMRDDBUS[9]);
buf (BRAMISOCMRDDBUS_delay[10], BRAMISOCMRDDBUS[10]);
buf (BRAMISOCMRDDBUS_delay[11], BRAMISOCMRDDBUS[11]);
buf (BRAMISOCMRDDBUS_delay[12], BRAMISOCMRDDBUS[12]);
buf (BRAMISOCMRDDBUS_delay[13], BRAMISOCMRDDBUS[13]);
buf (BRAMISOCMRDDBUS_delay[14], BRAMISOCMRDDBUS[14]);
buf (BRAMISOCMRDDBUS_delay[15], BRAMISOCMRDDBUS[15]);
buf (BRAMISOCMRDDBUS_delay[16], BRAMISOCMRDDBUS[16]);
buf (BRAMISOCMRDDBUS_delay[17], BRAMISOCMRDDBUS[17]);
buf (BRAMISOCMRDDBUS_delay[18], BRAMISOCMRDDBUS[18]);
buf (BRAMISOCMRDDBUS_delay[19], BRAMISOCMRDDBUS[19]);
buf (BRAMISOCMRDDBUS_delay[20], BRAMISOCMRDDBUS[20]);
buf (BRAMISOCMRDDBUS_delay[21], BRAMISOCMRDDBUS[21]);
buf (BRAMISOCMRDDBUS_delay[22], BRAMISOCMRDDBUS[22]);
buf (BRAMISOCMRDDBUS_delay[23], BRAMISOCMRDDBUS[23]);
buf (BRAMISOCMRDDBUS_delay[24], BRAMISOCMRDDBUS[24]);
buf (BRAMISOCMRDDBUS_delay[25], BRAMISOCMRDDBUS[25]);
buf (BRAMISOCMRDDBUS_delay[26], BRAMISOCMRDDBUS[26]);
buf (BRAMISOCMRDDBUS_delay[27], BRAMISOCMRDDBUS[27]);
buf (BRAMISOCMRDDBUS_delay[28], BRAMISOCMRDDBUS[28]);
buf (BRAMISOCMRDDBUS_delay[29], BRAMISOCMRDDBUS[29]);
buf (BRAMISOCMRDDBUS_delay[30], BRAMISOCMRDDBUS[30]);
buf (BRAMISOCMRDDBUS_delay[31], BRAMISOCMRDDBUS[31]);
buf (BRAMISOCMRDDBUS_delay[32], BRAMISOCMRDDBUS[32]);
buf (BRAMISOCMRDDBUS_delay[33], BRAMISOCMRDDBUS[33]);
buf (BRAMISOCMRDDBUS_delay[34], BRAMISOCMRDDBUS[34]);
buf (BRAMISOCMRDDBUS_delay[35], BRAMISOCMRDDBUS[35]);
buf (BRAMISOCMRDDBUS_delay[36], BRAMISOCMRDDBUS[36]);
buf (BRAMISOCMRDDBUS_delay[37], BRAMISOCMRDDBUS[37]);
buf (BRAMISOCMRDDBUS_delay[38], BRAMISOCMRDDBUS[38]);
buf (BRAMISOCMRDDBUS_delay[39], BRAMISOCMRDDBUS[39]);
buf (BRAMISOCMRDDBUS_delay[40], BRAMISOCMRDDBUS[40]);
buf (BRAMISOCMRDDBUS_delay[41], BRAMISOCMRDDBUS[41]);
buf (BRAMISOCMRDDBUS_delay[42], BRAMISOCMRDDBUS[42]);
buf (BRAMISOCMRDDBUS_delay[43], BRAMISOCMRDDBUS[43]);
buf (BRAMISOCMRDDBUS_delay[44], BRAMISOCMRDDBUS[44]);
buf (BRAMISOCMRDDBUS_delay[45], BRAMISOCMRDDBUS[45]);
buf (BRAMISOCMRDDBUS_delay[46], BRAMISOCMRDDBUS[46]);
buf (BRAMISOCMRDDBUS_delay[47], BRAMISOCMRDDBUS[47]);
buf (BRAMISOCMRDDBUS_delay[48], BRAMISOCMRDDBUS[48]);
buf (BRAMISOCMRDDBUS_delay[49], BRAMISOCMRDDBUS[49]);
buf (BRAMISOCMRDDBUS_delay[50], BRAMISOCMRDDBUS[50]);
buf (BRAMISOCMRDDBUS_delay[51], BRAMISOCMRDDBUS[51]);
buf (BRAMISOCMRDDBUS_delay[52], BRAMISOCMRDDBUS[52]);
buf (BRAMISOCMRDDBUS_delay[53], BRAMISOCMRDDBUS[53]);
buf (BRAMISOCMRDDBUS_delay[54], BRAMISOCMRDDBUS[54]);
buf (BRAMISOCMRDDBUS_delay[55], BRAMISOCMRDDBUS[55]);
buf (BRAMISOCMRDDBUS_delay[56], BRAMISOCMRDDBUS[56]);
buf (BRAMISOCMRDDBUS_delay[57], BRAMISOCMRDDBUS[57]);
buf (BRAMISOCMRDDBUS_delay[58], BRAMISOCMRDDBUS[58]);
buf (BRAMISOCMRDDBUS_delay[59], BRAMISOCMRDDBUS[59]);
buf (BRAMISOCMRDDBUS_delay[60], BRAMISOCMRDDBUS[60]);
buf (BRAMISOCMRDDBUS_delay[61], BRAMISOCMRDDBUS[61]);
buf (BRAMISOCMRDDBUS_delay[62], BRAMISOCMRDDBUS[62]);
buf (BRAMISOCMRDDBUS_delay[63], BRAMISOCMRDDBUS[63]);
buf (CPMC405CLOCK_delay, CPMC405CLOCK);
buf (CPMC405CORECLKINACTIVE_delay, CPMC405CORECLKINACTIVE);
buf (CPMC405CPUCLKEN_delay, CPMC405CPUCLKEN);
buf (CPMC405JTAGCLKEN_delay, CPMC405JTAGCLKEN);
buf (CPMC405TIMERCLKEN_delay, CPMC405TIMERCLKEN);
buf (CPMC405TIMERTICK_delay, CPMC405TIMERTICK);
buf (DBGC405DEBUGHALT_delay, DBGC405DEBUGHALT);
buf (DBGC405EXTBUSHOLDACK_delay, DBGC405EXTBUSHOLDACK);
buf (DBGC405UNCONDDEBUGEVENT_delay, DBGC405UNCONDDEBUGEVENT);
buf (DCRC405ACK_delay, DCRC405ACK);
buf (DCRC405DBUSIN_delay[0], DCRC405DBUSIN[0]);
buf (DCRC405DBUSIN_delay[1], DCRC405DBUSIN[1]);
buf (DCRC405DBUSIN_delay[2], DCRC405DBUSIN[2]);
buf (DCRC405DBUSIN_delay[3], DCRC405DBUSIN[3]);
buf (DCRC405DBUSIN_delay[4], DCRC405DBUSIN[4]);
buf (DCRC405DBUSIN_delay[5], DCRC405DBUSIN[5]);
buf (DCRC405DBUSIN_delay[6], DCRC405DBUSIN[6]);
buf (DCRC405DBUSIN_delay[7], DCRC405DBUSIN[7]);
buf (DCRC405DBUSIN_delay[8], DCRC405DBUSIN[8]);
buf (DCRC405DBUSIN_delay[9], DCRC405DBUSIN[9]);
buf (DCRC405DBUSIN_delay[10], DCRC405DBUSIN[10]);
buf (DCRC405DBUSIN_delay[11], DCRC405DBUSIN[11]);
buf (DCRC405DBUSIN_delay[12], DCRC405DBUSIN[12]);
buf (DCRC405DBUSIN_delay[13], DCRC405DBUSIN[13]);
buf (DCRC405DBUSIN_delay[14], DCRC405DBUSIN[14]);
buf (DCRC405DBUSIN_delay[15], DCRC405DBUSIN[15]);
buf (DCRC405DBUSIN_delay[16], DCRC405DBUSIN[16]);
buf (DCRC405DBUSIN_delay[17], DCRC405DBUSIN[17]);
buf (DCRC405DBUSIN_delay[18], DCRC405DBUSIN[18]);
buf (DCRC405DBUSIN_delay[19], DCRC405DBUSIN[19]);
buf (DCRC405DBUSIN_delay[20], DCRC405DBUSIN[20]);
buf (DCRC405DBUSIN_delay[21], DCRC405DBUSIN[21]);
buf (DCRC405DBUSIN_delay[22], DCRC405DBUSIN[22]);
buf (DCRC405DBUSIN_delay[23], DCRC405DBUSIN[23]);
buf (DCRC405DBUSIN_delay[24], DCRC405DBUSIN[24]);
buf (DCRC405DBUSIN_delay[25], DCRC405DBUSIN[25]);
buf (DCRC405DBUSIN_delay[26], DCRC405DBUSIN[26]);
buf (DCRC405DBUSIN_delay[27], DCRC405DBUSIN[27]);
buf (DCRC405DBUSIN_delay[28], DCRC405DBUSIN[28]);
buf (DCRC405DBUSIN_delay[29], DCRC405DBUSIN[29]);
buf (DCRC405DBUSIN_delay[30], DCRC405DBUSIN[30]);
buf (DCRC405DBUSIN_delay[31], DCRC405DBUSIN[31]);
buf (DSARCVALUE_delay[0], DSARCVALUE[0]);
buf (DSARCVALUE_delay[1], DSARCVALUE[1]);
buf (DSARCVALUE_delay[2], DSARCVALUE[2]);
buf (DSARCVALUE_delay[3], DSARCVALUE[3]);
buf (DSARCVALUE_delay[4], DSARCVALUE[4]);
buf (DSARCVALUE_delay[5], DSARCVALUE[5]);
buf (DSARCVALUE_delay[6], DSARCVALUE[6]);
buf (DSARCVALUE_delay[7], DSARCVALUE[7]);
buf (DSCNTLVALUE_delay[0], DSCNTLVALUE[0]);
buf (DSCNTLVALUE_delay[1], DSCNTLVALUE[1]);
buf (DSCNTLVALUE_delay[2], DSCNTLVALUE[2]);
buf (DSCNTLVALUE_delay[3], DSCNTLVALUE[3]);
buf (DSCNTLVALUE_delay[4], DSCNTLVALUE[4]);
buf (DSCNTLVALUE_delay[5], DSCNTLVALUE[5]);
buf (DSCNTLVALUE_delay[6], DSCNTLVALUE[6]);
buf (DSCNTLVALUE_delay[7], DSCNTLVALUE[7]);
buf (EICC405CRITINPUTIRQ_delay, EICC405CRITINPUTIRQ);
buf (EICC405EXTINPUTIRQ_delay, EICC405EXTINPUTIRQ);
// buf (GSR_delay, GSR);
buf (ISARCVALUE_delay[0], ISARCVALUE[0]);
buf (ISARCVALUE_delay[1], ISARCVALUE[1]);
buf (ISARCVALUE_delay[2], ISARCVALUE[2]);
buf (ISARCVALUE_delay[3], ISARCVALUE[3]);
buf (ISARCVALUE_delay[4], ISARCVALUE[4]);
buf (ISARCVALUE_delay[5], ISARCVALUE[5]);
buf (ISARCVALUE_delay[6], ISARCVALUE[6]);
buf (ISARCVALUE_delay[7], ISARCVALUE[7]);
buf (ISCNTLVALUE_delay[0], ISCNTLVALUE[0]);
buf (ISCNTLVALUE_delay[1], ISCNTLVALUE[1]);
buf (ISCNTLVALUE_delay[2], ISCNTLVALUE[2]);
buf (ISCNTLVALUE_delay[3], ISCNTLVALUE[3]);
buf (ISCNTLVALUE_delay[4], ISCNTLVALUE[4]);
buf (ISCNTLVALUE_delay[5], ISCNTLVALUE[5]);
buf (ISCNTLVALUE_delay[6], ISCNTLVALUE[6]);
buf (ISCNTLVALUE_delay[7], ISCNTLVALUE[7]);
buf (JTGC405BNDSCANTDO_delay, JTGC405BNDSCANTDO);
buf (JTGC405TCK_delay, JTGC405TCK);
buf (JTGC405TDI_delay, JTGC405TDI);
buf (JTGC405TMS_delay, JTGC405TMS);
buf (JTGC405TRSTNEG_delay, JTGC405TRSTNEG);
buf (MCBCPUCLKEN_delay, MCBCPUCLKEN);
buf (MCBJTAGEN_delay, MCBJTAGEN);
buf (MCBTIMEREN_delay, MCBTIMEREN);
buf (MCPPCRST_delay, MCPPCRST);
buf (PLBC405DCUADDRACK_delay, PLBC405DCUADDRACK);
buf (PLBC405DCUBUSY_delay, PLBC405DCUBUSY);
buf (PLBC405DCUERR_delay, PLBC405DCUERR);
buf (PLBC405DCURDDACK_delay, PLBC405DCURDDACK);
buf (PLBC405DCURDDBUS_delay[0], PLBC405DCURDDBUS[0]);
buf (PLBC405DCURDDBUS_delay[1], PLBC405DCURDDBUS[1]);
buf (PLBC405DCURDDBUS_delay[2], PLBC405DCURDDBUS[2]);
buf (PLBC405DCURDDBUS_delay[3], PLBC405DCURDDBUS[3]);
buf (PLBC405DCURDDBUS_delay[4], PLBC405DCURDDBUS[4]);
buf (PLBC405DCURDDBUS_delay[5], PLBC405DCURDDBUS[5]);
buf (PLBC405DCURDDBUS_delay[6], PLBC405DCURDDBUS[6]);
buf (PLBC405DCURDDBUS_delay[7], PLBC405DCURDDBUS[7]);
buf (PLBC405DCURDDBUS_delay[8], PLBC405DCURDDBUS[8]);
buf (PLBC405DCURDDBUS_delay[9], PLBC405DCURDDBUS[9]);
buf (PLBC405DCURDDBUS_delay[10], PLBC405DCURDDBUS[10]);
buf (PLBC405DCURDDBUS_delay[11], PLBC405DCURDDBUS[11]);
buf (PLBC405DCURDDBUS_delay[12], PLBC405DCURDDBUS[12]);
buf (PLBC405DCURDDBUS_delay[13], PLBC405DCURDDBUS[13]);
buf (PLBC405DCURDDBUS_delay[14], PLBC405DCURDDBUS[14]);
buf (PLBC405DCURDDBUS_delay[15], PLBC405DCURDDBUS[15]);
buf (PLBC405DCURDDBUS_delay[16], PLBC405DCURDDBUS[16]);
buf (PLBC405DCURDDBUS_delay[17], PLBC405DCURDDBUS[17]);
buf (PLBC405DCURDDBUS_delay[18], PLBC405DCURDDBUS[18]);
buf (PLBC405DCURDDBUS_delay[19], PLBC405DCURDDBUS[19]);
buf (PLBC405DCURDDBUS_delay[20], PLBC405DCURDDBUS[20]);
buf (PLBC405DCURDDBUS_delay[21], PLBC405DCURDDBUS[21]);
buf (PLBC405DCURDDBUS_delay[22], PLBC405DCURDDBUS[22]);
buf (PLBC405DCURDDBUS_delay[23], PLBC405DCURDDBUS[23]);
buf (PLBC405DCURDDBUS_delay[24], PLBC405DCURDDBUS[24]);
buf (PLBC405DCURDDBUS_delay[25], PLBC405DCURDDBUS[25]);
buf (PLBC405DCURDDBUS_delay[26], PLBC405DCURDDBUS[26]);
buf (PLBC405DCURDDBUS_delay[27], PLBC405DCURDDBUS[27]);
buf (PLBC405DCURDDBUS_delay[28], PLBC405DCURDDBUS[28]);
buf (PLBC405DCURDDBUS_delay[29], PLBC405DCURDDBUS[29]);
buf (PLBC405DCURDDBUS_delay[30], PLBC405DCURDDBUS[30]);
buf (PLBC405DCURDDBUS_delay[31], PLBC405DCURDDBUS[31]);
buf (PLBC405DCURDDBUS_delay[32], PLBC405DCURDDBUS[32]);
buf (PLBC405DCURDDBUS_delay[33], PLBC405DCURDDBUS[33]);
buf (PLBC405DCURDDBUS_delay[34], PLBC405DCURDDBUS[34]);
buf (PLBC405DCURDDBUS_delay[35], PLBC405DCURDDBUS[35]);
buf (PLBC405DCURDDBUS_delay[36], PLBC405DCURDDBUS[36]);
buf (PLBC405DCURDDBUS_delay[37], PLBC405DCURDDBUS[37]);
buf (PLBC405DCURDDBUS_delay[38], PLBC405DCURDDBUS[38]);
buf (PLBC405DCURDDBUS_delay[39], PLBC405DCURDDBUS[39]);
buf (PLBC405DCURDDBUS_delay[40], PLBC405DCURDDBUS[40]);
buf (PLBC405DCURDDBUS_delay[41], PLBC405DCURDDBUS[41]);
buf (PLBC405DCURDDBUS_delay[42], PLBC405DCURDDBUS[42]);
buf (PLBC405DCURDDBUS_delay[43], PLBC405DCURDDBUS[43]);
buf (PLBC405DCURDDBUS_delay[44], PLBC405DCURDDBUS[44]);
buf (PLBC405DCURDDBUS_delay[45], PLBC405DCURDDBUS[45]);
buf (PLBC405DCURDDBUS_delay[46], PLBC405DCURDDBUS[46]);
buf (PLBC405DCURDDBUS_delay[47], PLBC405DCURDDBUS[47]);
buf (PLBC405DCURDDBUS_delay[48], PLBC405DCURDDBUS[48]);
buf (PLBC405DCURDDBUS_delay[49], PLBC405DCURDDBUS[49]);
buf (PLBC405DCURDDBUS_delay[50], PLBC405DCURDDBUS[50]);
buf (PLBC405DCURDDBUS_delay[51], PLBC405DCURDDBUS[51]);
buf (PLBC405DCURDDBUS_delay[52], PLBC405DCURDDBUS[52]);
buf (PLBC405DCURDDBUS_delay[53], PLBC405DCURDDBUS[53]);
buf (PLBC405DCURDDBUS_delay[54], PLBC405DCURDDBUS[54]);
buf (PLBC405DCURDDBUS_delay[55], PLBC405DCURDDBUS[55]);
buf (PLBC405DCURDDBUS_delay[56], PLBC405DCURDDBUS[56]);
buf (PLBC405DCURDDBUS_delay[57], PLBC405DCURDDBUS[57]);
buf (PLBC405DCURDDBUS_delay[58], PLBC405DCURDDBUS[58]);
buf (PLBC405DCURDDBUS_delay[59], PLBC405DCURDDBUS[59]);
buf (PLBC405DCURDDBUS_delay[60], PLBC405DCURDDBUS[60]);
buf (PLBC405DCURDDBUS_delay[61], PLBC405DCURDDBUS[61]);
buf (PLBC405DCURDDBUS_delay[62], PLBC405DCURDDBUS[62]);
buf (PLBC405DCURDDBUS_delay[63], PLBC405DCURDDBUS[63]);
buf (PLBC405DCURDWDADDR_delay[1], PLBC405DCURDWDADDR[1]);
buf (PLBC405DCURDWDADDR_delay[2], PLBC405DCURDWDADDR[2]);
buf (PLBC405DCURDWDADDR_delay[3], PLBC405DCURDWDADDR[3]);
buf (PLBC405DCUSSIZE1_delay, PLBC405DCUSSIZE1);
buf (PLBC405DCUWRDACK_delay, PLBC405DCUWRDACK);
buf (PLBC405ICUADDRACK_delay, PLBC405ICUADDRACK);
buf (PLBC405ICUBUSY_delay, PLBC405ICUBUSY);
buf (PLBC405ICUERR_delay, PLBC405ICUERR);
buf (PLBC405ICURDDACK_delay, PLBC405ICURDDACK);
buf (PLBC405ICURDDBUS_delay[0], PLBC405ICURDDBUS[0]);
buf (PLBC405ICURDDBUS_delay[1], PLBC405ICURDDBUS[1]);
buf (PLBC405ICURDDBUS_delay[2], PLBC405ICURDDBUS[2]);
buf (PLBC405ICURDDBUS_delay[3], PLBC405ICURDDBUS[3]);
buf (PLBC405ICURDDBUS_delay[4], PLBC405ICURDDBUS[4]);
buf (PLBC405ICURDDBUS_delay[5], PLBC405ICURDDBUS[5]);
buf (PLBC405ICURDDBUS_delay[6], PLBC405ICURDDBUS[6]);
buf (PLBC405ICURDDBUS_delay[7], PLBC405ICURDDBUS[7]);
buf (PLBC405ICURDDBUS_delay[8], PLBC405ICURDDBUS[8]);
buf (PLBC405ICURDDBUS_delay[9], PLBC405ICURDDBUS[9]);
buf (PLBC405ICURDDBUS_delay[10], PLBC405ICURDDBUS[10]);
buf (PLBC405ICURDDBUS_delay[11], PLBC405ICURDDBUS[11]);
buf (PLBC405ICURDDBUS_delay[12], PLBC405ICURDDBUS[12]);
buf (PLBC405ICURDDBUS_delay[13], PLBC405ICURDDBUS[13]);
buf (PLBC405ICURDDBUS_delay[14], PLBC405ICURDDBUS[14]);
buf (PLBC405ICURDDBUS_delay[15], PLBC405ICURDDBUS[15]);
buf (PLBC405ICURDDBUS_delay[16], PLBC405ICURDDBUS[16]);
buf (PLBC405ICURDDBUS_delay[17], PLBC405ICURDDBUS[17]);
buf (PLBC405ICURDDBUS_delay[18], PLBC405ICURDDBUS[18]);
buf (PLBC405ICURDDBUS_delay[19], PLBC405ICURDDBUS[19]);
buf (PLBC405ICURDDBUS_delay[20], PLBC405ICURDDBUS[20]);
buf (PLBC405ICURDDBUS_delay[21], PLBC405ICURDDBUS[21]);
buf (PLBC405ICURDDBUS_delay[22], PLBC405ICURDDBUS[22]);
buf (PLBC405ICURDDBUS_delay[23], PLBC405ICURDDBUS[23]);
buf (PLBC405ICURDDBUS_delay[24], PLBC405ICURDDBUS[24]);
buf (PLBC405ICURDDBUS_delay[25], PLBC405ICURDDBUS[25]);
buf (PLBC405ICURDDBUS_delay[26], PLBC405ICURDDBUS[26]);
buf (PLBC405ICURDDBUS_delay[27], PLBC405ICURDDBUS[27]);
buf (PLBC405ICURDDBUS_delay[28], PLBC405ICURDDBUS[28]);
buf (PLBC405ICURDDBUS_delay[29], PLBC405ICURDDBUS[29]);
buf (PLBC405ICURDDBUS_delay[30], PLBC405ICURDDBUS[30]);
buf (PLBC405ICURDDBUS_delay[31], PLBC405ICURDDBUS[31]);
buf (PLBC405ICURDDBUS_delay[32], PLBC405ICURDDBUS[32]);
buf (PLBC405ICURDDBUS_delay[33], PLBC405ICURDDBUS[33]);
buf (PLBC405ICURDDBUS_delay[34], PLBC405ICURDDBUS[34]);
buf (PLBC405ICURDDBUS_delay[35], PLBC405ICURDDBUS[35]);
buf (PLBC405ICURDDBUS_delay[36], PLBC405ICURDDBUS[36]);
buf (PLBC405ICURDDBUS_delay[37], PLBC405ICURDDBUS[37]);
buf (PLBC405ICURDDBUS_delay[38], PLBC405ICURDDBUS[38]);
buf (PLBC405ICURDDBUS_delay[39], PLBC405ICURDDBUS[39]);
buf (PLBC405ICURDDBUS_delay[40], PLBC405ICURDDBUS[40]);
buf (PLBC405ICURDDBUS_delay[41], PLBC405ICURDDBUS[41]);
buf (PLBC405ICURDDBUS_delay[42], PLBC405ICURDDBUS[42]);
buf (PLBC405ICURDDBUS_delay[43], PLBC405ICURDDBUS[43]);
buf (PLBC405ICURDDBUS_delay[44], PLBC405ICURDDBUS[44]);
buf (PLBC405ICURDDBUS_delay[45], PLBC405ICURDDBUS[45]);
buf (PLBC405ICURDDBUS_delay[46], PLBC405ICURDDBUS[46]);
buf (PLBC405ICURDDBUS_delay[47], PLBC405ICURDDBUS[47]);
buf (PLBC405ICURDDBUS_delay[48], PLBC405ICURDDBUS[48]);
buf (PLBC405ICURDDBUS_delay[49], PLBC405ICURDDBUS[49]);
buf (PLBC405ICURDDBUS_delay[50], PLBC405ICURDDBUS[50]);
buf (PLBC405ICURDDBUS_delay[51], PLBC405ICURDDBUS[51]);
buf (PLBC405ICURDDBUS_delay[52], PLBC405ICURDDBUS[52]);
buf (PLBC405ICURDDBUS_delay[53], PLBC405ICURDDBUS[53]);
buf (PLBC405ICURDDBUS_delay[54], PLBC405ICURDDBUS[54]);
buf (PLBC405ICURDDBUS_delay[55], PLBC405ICURDDBUS[55]);
buf (PLBC405ICURDDBUS_delay[56], PLBC405ICURDDBUS[56]);
buf (PLBC405ICURDDBUS_delay[57], PLBC405ICURDDBUS[57]);
buf (PLBC405ICURDDBUS_delay[58], PLBC405ICURDDBUS[58]);
buf (PLBC405ICURDDBUS_delay[59], PLBC405ICURDDBUS[59]);
buf (PLBC405ICURDDBUS_delay[60], PLBC405ICURDDBUS[60]);
buf (PLBC405ICURDDBUS_delay[61], PLBC405ICURDDBUS[61]);
buf (PLBC405ICURDDBUS_delay[62], PLBC405ICURDDBUS[62]);
buf (PLBC405ICURDDBUS_delay[63], PLBC405ICURDDBUS[63]);
buf (PLBC405ICURDWDADDR_delay[1], PLBC405ICURDWDADDR[1]);
buf (PLBC405ICURDWDADDR_delay[2], PLBC405ICURDWDADDR[2]);
buf (PLBC405ICURDWDADDR_delay[3], PLBC405ICURDWDADDR[3]);
buf (PLBC405ICUSSIZE1_delay, PLBC405ICUSSIZE1);
buf (PLBCLK_delay, PLBCLK);
buf (RSTC405RESETCHIP_delay, RSTC405RESETCHIP);
buf (RSTC405RESETCORE_delay, RSTC405RESETCORE);
buf (RSTC405RESETSYS_delay, RSTC405RESETSYS);
buf (TIEC405DETERMINISTICMULT_delay, TIEC405DETERMINISTICMULT);
buf (TIEC405DISOPERANDFWD_delay, TIEC405DISOPERANDFWD);
buf (TIEC405MMUEN_delay, TIEC405MMUEN);
buf (TIEDSOCMDCRADDR_delay[0], TIEDSOCMDCRADDR[0]);
buf (TIEDSOCMDCRADDR_delay[1], TIEDSOCMDCRADDR[1]);
buf (TIEDSOCMDCRADDR_delay[2], TIEDSOCMDCRADDR[2]);
buf (TIEDSOCMDCRADDR_delay[3], TIEDSOCMDCRADDR[3]);
buf (TIEDSOCMDCRADDR_delay[4], TIEDSOCMDCRADDR[4]);
buf (TIEDSOCMDCRADDR_delay[5], TIEDSOCMDCRADDR[5]);
buf (TIEDSOCMDCRADDR_delay[6], TIEDSOCMDCRADDR[6]);
buf (TIEDSOCMDCRADDR_delay[7], TIEDSOCMDCRADDR[7]);
buf (TIEISOCMDCRADDR_delay[0], TIEISOCMDCRADDR[0]);
buf (TIEISOCMDCRADDR_delay[1], TIEISOCMDCRADDR[1]);
buf (TIEISOCMDCRADDR_delay[2], TIEISOCMDCRADDR[2]);
buf (TIEISOCMDCRADDR_delay[3], TIEISOCMDCRADDR[3]);
buf (TIEISOCMDCRADDR_delay[4], TIEISOCMDCRADDR[4]);
buf (TIEISOCMDCRADDR_delay[5], TIEISOCMDCRADDR[5]);
buf (TIEISOCMDCRADDR_delay[6], TIEISOCMDCRADDR[6]);
buf (TIEISOCMDCRADDR_delay[7], TIEISOCMDCRADDR[7]);
buf (TRCC405TRACEDISABLE_delay, TRCC405TRACEDISABLE);
buf (TRCC405TRIGGEREVENTIN_delay, TRCC405TRIGGEREVENTIN);

wire    FPGA_CCLK;
wire	FPGA_BUS_RESET;
wire	FPGA_GSR;
wire	FPGA_GWE;
wire	FPGA_GHIGHB;
wire	GSR_OR;

reg	FPGA_POR;
reg	FPGA_CCLK_REG;

`ifdef STARTUP_BLK
	assign FPGA_CCLK	= TESTBENCH.FPGA_cclk;
	assign  FPGA_BUS_RESET 	= TESTBENCH.FPGA_bus_reset;
	assign  GSR_OR 		= TESTBENCH.FPGA_gsr;
	assign  FPGA_GWE 	= TESTBENCH.FPGA_gwe;
	assign  FPGA_GHIGHB 	= TESTBENCH.FPGA_ghigh_b;
`else

FPGA_startup start_blk(
.bus_reset	(FPGA_BUS_RESET),
.ghigh_b	(FPGA_GHIGHB), 
.gsr		(FPGA_GSR), 
.done		(), 
.gwe		(FPGA_GWE), 
.gts_b		(), 
.shutdown	(1'b0), 
.cclk		(FPGA_CCLK), 
.por		(FPGA_POR)
);

or IGSR_OR (GSR_OR, FPGA_GSR, GSR);

`define Loc_FPGA_POR_TIME           10   // FPGA Power-On Reset time

// Generate FPGA CCLK
 always
    #500 FPGA_CCLK_REG = ~FPGA_CCLK_REG;

assign FPGA_CCLK = FPGA_CCLK_REG;

initial begin
    FPGA_CCLK_REG = 0;
    FPGA_POR  = 1'b1;
    #(`Loc_FPGA_POR_TIME)       FPGA_POR  = 1'b0;
end

`endif   // STARTUP_BLK

wire FPGA_BUS_RESET_delay;
wire GSR_delay;
wire FPGA_GWE_delay;
wire FPGA_GHIGHB_delay;

assign #(in_delay) FPGA_BUS_RESET_delay = FPGA_BUS_RESET;
assign #(in_delay) GSR_delay = GSR_OR;
assign #(in_delay) FPGA_GWE_delay = FPGA_GWE;
assign #(in_delay) FPGA_GHIGHB_delay = FPGA_GHIGHB;

`ifdef ProcBlk_RTL
usr_proc_block_cap Iusr_proc_block_cap(
`else
PPC405_SWIFT IPPC405_SWIFT(
`endif          //ProcBlk_rtl

   .BUS_CLK(FPGA_CCLK),
   .BUS_RESET(FPGA_BUS_RESET_delay),
   .GSR(GSR_delay),
   .GWE(FPGA_GWE_delay),
   .GHIGHB(FPGA_GHIGHB_delay),
   .CPMC405CPUCLKEN(CPMC405CPUCLKEN_delay),
   .CPMC405JTAGCLKEN(CPMC405JTAGCLKEN_delay),
   .CPMC405TIMERCLKEN(CPMC405TIMERCLKEN_delay),
   .C405JTGPGMOUT(C405JTGPGMOUT_delay),
   .MCBCPUCLKEN(MCBCPUCLKEN_delay),
   .MCBJTAGEN(MCBJTAGEN_delay),
   .MCBTIMEREN(MCBTIMEREN_delay),
   .MCPPCRST(MCPPCRST_delay),
   .C405TRCODDEXECUTIONSTATUS(C405TRCODDEXECUTIONSTATUS_delay),
   .C405TRCEVENEXECUTIONSTATUS(C405TRCEVENEXECUTIONSTATUS_delay),
   .CPMC405CLOCK(CPMC405CLOCK_delay),
   .CPMC405CORECLKINACTIVE(CPMC405CORECLKINACTIVE_delay),
   .PLBCLK(PLBCLK_delay),
   .CPMC405TIMERTICK(CPMC405TIMERTICK_delay),
   .C405CPMMSREE(C405CPMMSREE_delay),
   .C405CPMMSRCE(C405CPMMSRCE_delay),
   .C405CPMTIMERIRQ(C405CPMTIMERIRQ_delay),
   .C405CPMTIMERRESETREQ(C405CPMTIMERRESETREQ_delay),
   .C405CPMCORESLEEPREQ(C405CPMCORESLEEPREQ_delay),
   .TIEC405DISOPERANDFWD(TIEC405DISOPERANDFWD_delay),
   .TIEC405DETERMINISTICMULT(TIEC405DETERMINISTICMULT_delay),
   .TIEC405MMUEN(TIEC405MMUEN_delay),
   .TIEC405PVR(PPCUSER),
   .C405XXXMACHINECHECK(C405XXXMACHINECHECK_delay),
   .C405RSTCHIPRESETREQ(C405RSTCHIPRESETREQ_delay),
   .C405RSTCORERESETREQ(C405RSTCORERESETREQ_delay),
   .C405RSTSYSRESETREQ(C405RSTSYSRESETREQ_delay),
   .RSTC405RESETCHIP(RSTC405RESETCHIP_delay),
   .RSTC405RESETCORE(RSTC405RESETCORE_delay),
   .RSTC405RESETSYS(RSTC405RESETSYS_delay),
   .C405PLBICUREQUEST(C405PLBICUREQUEST_delay),
   .C405PLBICUPRIORITY(C405PLBICUPRIORITY_delay),
   .C405PLBICUCACHEABLE(C405PLBICUCACHEABLE_delay),
   .C405PLBICUABUS(C405PLBICUABUS_delay),
   .C405PLBICUSIZE(C405PLBICUSIZE_delay),
   .C405PLBICUABORT(C405PLBICUABORT_delay),
   .C405PLBICUU0ATTR(C405PLBICUU0ATTR_delay),
   .PLBC405ICUADDRACK(PLBC405ICUADDRACK_delay),
   .PLBC405ICUBUSY(PLBC405ICUBUSY_delay),
   .PLBC405ICUERR(PLBC405ICUERR_delay),
   .PLBC405ICURDDACK(PLBC405ICURDDACK_delay),
   .PLBC405ICURDDBUS(PLBC405ICURDDBUS_delay),
   .PLBC405ICUSSIZE1(PLBC405ICUSSIZE1_delay),
   .PLBC405ICURDWDADDR(PLBC405ICURDWDADDR_delay),
   .C405PLBDCUREQUEST(C405PLBDCUREQUEST_delay),
   .C405PLBDCURNW(C405PLBDCURNW_delay),
   .C405PLBDCUABUS(C405PLBDCUABUS_delay),
   .C405PLBDCUBE(C405PLBDCUBE_delay),
   .C405PLBDCUCACHEABLE(C405PLBDCUCACHEABLE_delay),
   .C405PLBDCUGUARDED(C405PLBDCUGUARDED_delay),
   .C405PLBDCUPRIORITY(C405PLBDCUPRIORITY_delay),
   .C405PLBDCUSIZE2(C405PLBDCUSIZE2_delay),
   .C405PLBDCUABORT(C405PLBDCUABORT_delay),
   .C405PLBDCUWRDBUS(C405PLBDCUWRDBUS_delay),
   .C405PLBDCUU0ATTR(C405PLBDCUU0ATTR_delay),
   .C405PLBDCUWRITETHRU(C405PLBDCUWRITETHRU_delay),
   .PLBC405DCUADDRACK(PLBC405DCUADDRACK_delay),
   .PLBC405DCUBUSY(PLBC405DCUBUSY_delay),
   .PLBC405DCUERR(PLBC405DCUERR_delay),
   .PLBC405DCURDDACK(PLBC405DCURDDACK_delay),
   .PLBC405DCURDDBUS(PLBC405DCURDDBUS_delay),
   .PLBC405DCURDWDADDR(PLBC405DCURDWDADDR_delay),
   .PLBC405DCUSSIZE1(PLBC405DCUSSIZE1_delay),
   .PLBC405DCUWRDACK(PLBC405DCUWRDACK_delay),
   .ISOCMBRAMRDABUS(ISOCMBRAMRDABUS_delay),
   .ISOCMBRAMWRABUS(ISOCMBRAMWRABUS_delay),
   .ISOCMBRAMEN(ISOCMBRAMEN_delay),
   .ISOCMBRAMODDWRITEEN(ISOCMBRAMODDWRITEEN_delay),
   .ISOCMBRAMEVENWRITEEN(ISOCMBRAMEVENWRITEEN_delay),
   .ISOCMBRAMWRDBUS(ISOCMBRAMWRDBUS_delay),
   .BRAMISOCMRDDBUS(BRAMISOCMRDDBUS_delay),
   .TIEISOCMDCRADDR(TIEISOCMDCRADDR_delay),
   .ISARCVALUE(ISARCVALUE_delay),
   .ISCNTLVALUE(ISCNTLVALUE_delay),
   .BRAMISOCMCLK(BRAMISOCMCLK_delay),
   .DSOCMBRAMABUS(DSOCMBRAMABUS_delay),
   .DSOCMBRAMBYTEWRITE(DSOCMBRAMBYTEWRITE_delay),
   .DSOCMBRAMEN(DSOCMBRAMEN_delay),
   .DSOCMBRAMWRDBUS(DSOCMBRAMWRDBUS_delay),
   .BRAMDSOCMRDDBUS(BRAMDSOCMRDDBUS_delay),
   .DSOCMBUSY(DSOCMBUSY_delay),
   .TIEDSOCMDCRADDR(TIEDSOCMDCRADDR_delay),
   .DSARCVALUE(DSARCVALUE_delay),
   .DSCNTLVALUE(DSCNTLVALUE_delay),
   .BRAMDSOCMCLK(BRAMDSOCMCLK_delay),
   .C405DCRREAD(C405DCRREAD_delay),
   .C405DCRWRITE(C405DCRWRITE_delay),
   .C405DCRABUS(C405DCRABUS_delay),
   .C405DCRDBUSOUT(C405DCRDBUSOUT_delay),
   .DCRC405ACK(DCRC405ACK_delay),
   .DCRC405DBUSIN(DCRC405DBUSIN_delay),
   .EICC405EXTINPUTIRQ(EICC405EXTINPUTIRQ_delay),
   .EICC405CRITINPUTIRQ(EICC405CRITINPUTIRQ_delay),
   .JTGC405BNDSCANTDO(JTGC405BNDSCANTDO_delay),
   .JTGC405TCK(JTGC405TCK_delay),
   .JTGC405TDI(JTGC405TDI_delay),
   .JTGC405TMS(JTGC405TMS_delay),
   .JTGC405TRSTNEG(JTGC405TRSTNEG_delay),
   .C405JTGTDO(C405JTGTDO_delay),
   .C405JTGTDOEN(C405JTGTDOEN_delay),
   .C405JTGEXTEST(C405JTGEXTEST_delay),
   .C405JTGCAPTUREDR(C405JTGCAPTUREDR_delay),
   .C405JTGSHIFTDR(C405JTGSHIFTDR_delay),
   .C405JTGUPDATEDR(C405JTGUPDATEDR_delay),
   .DBGC405DEBUGHALT(DBGC405DEBUGHALT_delay),
   .DBGC405UNCONDDEBUGEVENT(DBGC405UNCONDDEBUGEVENT_delay),
   .DBGC405EXTBUSHOLDACK(DBGC405EXTBUSHOLDACK_delay),
   .C405DBGMSRWE(C405DBGMSRWE_delay),
   .C405DBGSTOPACK(C405DBGSTOPACK_delay),
   .C405DBGWBCOMPLETE(C405DBGWBCOMPLETE_delay),
   .C405DBGWBFULL(C405DBGWBFULL_delay),
   .C405DBGWBIAR(C405DBGWBIAR_delay),
   .C405TRCTRIGGEREVENTOUT(C405TRCTRIGGEREVENTOUT_delay),
   .C405TRCTRIGGEREVENTTYPE(C405TRCTRIGGEREVENTTYPE_delay),
   .C405TRCCYCLE(C405TRCCYCLE_delay),
   .C405TRCTRACESTATUS(C405TRCTRACESTATUS_delay),
   .TRCC405TRACEDISABLE(TRCC405TRACEDISABLE_delay),
   .TRCC405TRIGGEREVENTIN(TRCC405TRIGGEREVENTIN_delay)
);

specify

	(BRAMISOCMCLK => ISOCMBRAMEN) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMEVENWRITEEN) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMODDWRITEEN) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[8]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[9]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[10]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[11]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[12]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[13]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[14]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[15]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[16]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[17]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[18]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[19]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[20]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[21]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[22]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[23]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[24]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[25]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[26]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[27]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMRDABUS[28]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[8]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[9]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[10]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[11]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[12]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[13]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[14]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[15]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[16]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[17]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[18]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[19]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[20]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[21]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[22]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[23]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[24]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[25]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[26]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[27]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRABUS[28]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[0]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[1]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[2]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[3]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[4]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[5]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[6]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[7]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[8]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[9]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[10]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[11]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[12]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[13]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[14]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[15]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[16]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[17]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[18]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[19]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[20]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[21]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[22]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[23]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[24]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[25]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[26]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[27]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[28]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[29]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[30]) = (0:0:0, 0:0:0);
	(BRAMISOCMCLK => ISOCMBRAMWRDBUS[31]) = (0:0:0, 0:0:0);

	(BRAMDSOCMCLK => DSOCMBRAMABUS[8]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[9]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[10]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[11]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[12]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[13]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[14]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[15]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[16]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[17]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[18]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[19]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[20]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[21]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[22]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[23]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[24]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[25]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[26]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[27]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[28]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMABUS[29]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMBYTEWRITE[0]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMBYTEWRITE[1]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMBYTEWRITE[2]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMBYTEWRITE[3]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMEN) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[0]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[1]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[2]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[3]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[4]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[5]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[6]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[7]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[8]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[9]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[10]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[11]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[12]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[13]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[14]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[15]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[16]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[17]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[18]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[19]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[20]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[21]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[22]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[23]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[24]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[25]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[26]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[27]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[28]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[29]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[30]) = (0:0:0, 0:0:0);
	(BRAMDSOCMCLK => DSOCMBRAMWRDBUS[31]) = (0:0:0, 0:0:0);

	(CPMC405CLOCK => C405CPMCORESLEEPREQ) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405CPMMSRCE) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405CPMMSREE) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405CPMTIMERIRQ) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405CPMTIMERRESETREQ) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGMSRWE) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGSTOPACK) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBCOMPLETE) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBFULL) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[2]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[3]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[4]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[5]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[6]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[7]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[8]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[9]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[10]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[11]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[12]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[13]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[14]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[15]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[16]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[17]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[18]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[19]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[20]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[21]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[22]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[23]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[24]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[25]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[26]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[27]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[28]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DBGWBIAR[29]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[2]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[3]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[4]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[5]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[6]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[7]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[8]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRABUS[9]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[2]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[3]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[4]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[5]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[6]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[7]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[8]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[9]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[10]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[11]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[12]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[13]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[14]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[15]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[16]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[17]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[18]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[19]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[20]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[21]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[22]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[23]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[24]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[25]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[26]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[27]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[28]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[29]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[30]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRDBUSOUT[31]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRREAD) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405DCRWRITE) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405JTGPGMOUT) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405RSTCHIPRESETREQ) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405RSTCORERESETREQ) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405RSTSYSRESETREQ) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCCYCLE) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCEVENEXECUTIONSTATUS[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCEVENEXECUTIONSTATUS[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCODDEXECUTIONSTATUS[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCODDEXECUTIONSTATUS[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRACESTATUS[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRACESTATUS[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRACESTATUS[2]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRACESTATUS[3]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTOUT) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[0]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[1]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[2]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[3]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[4]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[5]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[6]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[7]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[8]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[9]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405TRCTRIGGEREVENTTYPE[10]) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => C405XXXMACHINECHECK) = (0:0:0, 0:0:0);
	(CPMC405CLOCK => DSOCMBUSY) = (0:0:0, 0:0:0);

	(GSR => C405RSTCORERESETREQ) = (0:0:0, 0:0:0);

	(JTGC405TCK => C405JTGCAPTUREDR) = (0:0:0, 0:0:0);
	(JTGC405TCK => C405JTGEXTEST) = (0:0:0, 0:0:0);
	(JTGC405TCK => C405JTGSHIFTDR) = (0:0:0, 0:0:0);
	(JTGC405TCK => C405JTGTDO) = (0:0:0, 0:0:0);
	(JTGC405TCK => C405JTGTDOEN) = (0:0:0, 0:0:0);
	(JTGC405TCK => C405JTGUPDATEDR) = (0:0:0, 0:0:0);

	(PLBCLK => C405PLBDCUABORT) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[0]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[1]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[2]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[3]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[4]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[5]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[6]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[7]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[8]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[9]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[10]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[11]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[12]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[13]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[14]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[15]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[16]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[17]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[18]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[19]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[20]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[21]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[22]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[23]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[24]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[25]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[26]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[27]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[28]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[29]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[30]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUABUS[31]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[0]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[1]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[2]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[3]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[4]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[5]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[6]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUBE[7]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUCACHEABLE) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUGUARDED) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUPRIORITY[0]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUPRIORITY[1]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUREQUEST) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCURNW) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUSIZE2) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUU0ATTR) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[0]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[1]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[2]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[3]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[4]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[5]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[6]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[7]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[8]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[9]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[10]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[11]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[12]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[13]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[14]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[15]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[16]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[17]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[18]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[19]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[20]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[21]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[22]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[23]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[24]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[25]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[26]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[27]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[28]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[29]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[30]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[31]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[32]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[33]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[34]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[35]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[36]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[37]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[38]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[39]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[40]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[41]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[42]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[43]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[44]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[45]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[46]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[47]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[48]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[49]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[50]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[51]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[52]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[53]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[54]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[55]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[56]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[57]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[58]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[59]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[60]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[61]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[62]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRDBUS[63]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBDCUWRITETHRU) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABORT) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[0]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[1]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[2]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[3]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[4]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[5]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[6]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[7]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[8]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[9]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[10]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[11]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[12]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[13]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[14]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[15]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[16]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[17]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[18]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[19]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[20]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[21]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[22]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[23]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[24]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[25]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[26]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[27]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[28]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUABUS[29]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUCACHEABLE) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUPRIORITY[0]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUPRIORITY[1]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUREQUEST) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUSIZE[2]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUSIZE[3]) = (0:0:0, 0:0:0);
	(PLBCLK => C405PLBICUU0ATTR) = (0:0:0, 0:0:0);

	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, posedge BRAMDSOCMRDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMDSOCMCLK, negedge BRAMDSOCMRDDBUS[31], 0:0:0, 0:0:0);

	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[32], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[32], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[33], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[33], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[34], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[34], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[35], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[35], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[36], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[36], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[37], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[37], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[38], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[38], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[39], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[39], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[40], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[40], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[41], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[41], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[42], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[42], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[43], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[43], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[44], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[44], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[45], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[45], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[46], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[46], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[47], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[47], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[48], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[48], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[49], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[49], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[50], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[50], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[51], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[51], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[52], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[52], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[53], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[53], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[54], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[54], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[55], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[55], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[56], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[56], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[57], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[57], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[58], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[58], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[59], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[59], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[60], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[60], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[61], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[61], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[62], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[62], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, posedge BRAMISOCMRDDBUS[63], 0:0:0, 0:0:0);
	$setuphold (posedge BRAMISOCMCLK, negedge BRAMISOCMRDDBUS[63], 0:0:0, 0:0:0);

	$setuphold (posedge CPMC405CLOCK, posedge CPMC405CPUCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge CPMC405CPUCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge CPMC405JTAGCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge CPMC405JTAGCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge CPMC405TIMERCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge CPMC405TIMERCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge CPMC405TIMERTICK, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge CPMC405TIMERTICK, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DBGC405DEBUGHALT, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DBGC405DEBUGHALT, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DBGC405UNCONDDEBUGEVENT, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DBGC405UNCONDDEBUGEVENT, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405ACK, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405ACK, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[8], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[8], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[9], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[9], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[10], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[10], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[11], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[11], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[12], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[12], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[13], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[13], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[14], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[14], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[15], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[15], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[16], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[16], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[17], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[17], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[18], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[18], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[19], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[19], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[20], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[20], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[21], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[21], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[22], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[22], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[23], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[23], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[24], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[24], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[25], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[25], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[26], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[26], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[27], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[27], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[28], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[28], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[29], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[29], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[30], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[30], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DCRC405DBUSIN[31], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DCRC405DBUSIN[31], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSARCVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSARCVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge DSCNTLVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge DSCNTLVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge EICC405CRITINPUTIRQ, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge EICC405CRITINPUTIRQ, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge EICC405EXTINPUTIRQ, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge EICC405EXTINPUTIRQ, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISARCVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISARCVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge ISCNTLVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge ISCNTLVALUE[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge MCBCPUCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge MCBCPUCLKEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge MCBJTAGEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge MCBJTAGEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge MCBTIMEREN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge MCBTIMEREN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge MCPPCRST, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge MCPPCRST, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge PLBCLK, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge PLBCLK, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge RSTC405RESETCHIP, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge RSTC405RESETCHIP, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge RSTC405RESETCORE, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge RSTC405RESETCORE, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge RSTC405RESETSYS, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge RSTC405RESETSYS, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEC405DETERMINISTICMULT, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEC405DETERMINISTICMULT, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEC405DISOPERANDFWD, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEC405DISOPERANDFWD, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEC405MMUEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEC405MMUEN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEDSOCMDCRADDR[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEDSOCMDCRADDR[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[0], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[4], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[5], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[6], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TIEISOCMDCRADDR[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TIEISOCMDCRADDR[7], 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TRCC405TRACEDISABLE, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TRCC405TRACEDISABLE, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, posedge TRCC405TRIGGEREVENTIN, 0:0:0, 0:0:0);
	$setuphold (posedge CPMC405CLOCK, negedge TRCC405TRIGGEREVENTIN, 0:0:0, 0:0:0);

	$setuphold (posedge JTGC405TCK, posedge CPMC405CORECLKINACTIVE, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, negedge CPMC405CORECLKINACTIVE, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, posedge DBGC405EXTBUSHOLDACK, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, negedge DBGC405EXTBUSHOLDACK, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, posedge JTGC405BNDSCANTDO, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, negedge JTGC405BNDSCANTDO, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, posedge JTGC405TDI, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, negedge JTGC405TDI, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, posedge JTGC405TMS, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, negedge JTGC405TMS, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, posedge JTGC405TRSTNEG, 0:0:0, 0:0:0);
	$setuphold (posedge JTGC405TCK, negedge JTGC405TRSTNEG, 0:0:0, 0:0:0);

	$setuphold (posedge PLBCLK, posedge PLBC405DCUADDRACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCUADDRACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCUBUSY, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCUBUSY, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCUERR, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCUERR, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[32], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[32], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[33], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[33], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[34], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[34], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[35], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[35], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[36], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[36], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[37], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[37], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[38], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[38], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[39], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[39], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[40], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[40], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[41], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[41], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[42], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[42], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[43], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[43], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[44], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[44], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[45], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[45], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[46], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[46], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[47], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[47], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[48], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[48], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[49], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[49], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[50], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[50], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[51], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[51], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[52], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[52], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[53], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[53], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[54], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[54], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[55], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[55], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[56], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[56], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[57], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[57], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[58], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[58], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[59], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[59], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[60], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[60], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[61], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[61], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[62], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[62], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDDBUS[63], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDDBUS[63], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDWDADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDWDADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDWDADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDWDADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCURDWDADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCURDWDADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCUSSIZE1, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCUSSIZE1, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405DCUWRDACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405DCUWRDACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICUADDRACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICUADDRACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICUBUSY, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICUBUSY, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICUERR, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICUERR, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDACK, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[0], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[4], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[5], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[6], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[7], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[8], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[9], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[10], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[11], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[12], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[13], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[14], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[15], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[16], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[17], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[18], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[19], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[20], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[21], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[22], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[23], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[24], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[25], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[26], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[27], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[28], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[29], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[30], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[31], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[32], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[32], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[33], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[33], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[34], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[34], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[35], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[35], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[36], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[36], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[37], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[37], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[38], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[38], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[39], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[39], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[40], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[40], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[41], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[41], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[42], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[42], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[43], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[43], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[44], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[44], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[45], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[45], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[46], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[46], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[47], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[47], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[48], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[48], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[49], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[49], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[50], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[50], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[51], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[51], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[52], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[52], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[53], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[53], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[54], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[54], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[55], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[55], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[56], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[56], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[57], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[57], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[58], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[58], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[59], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[59], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[60], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[60], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[61], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[61], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[62], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[62], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDDBUS[63], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDDBUS[63], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDWDADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDWDADDR[1], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDWDADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDWDADDR[2], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICURDWDADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICURDWDADDR[3], 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, posedge PLBC405ICUSSIZE1, 0:0:0, 0:0:0);
	$setuphold (posedge PLBCLK, negedge PLBC405ICUSSIZE1, 0:0:0, 0:0:0);

	$width (posedge BRAMDSOCMCLK, 0:0:0, 0, notifier);
	$width (negedge BRAMDSOCMCLK, 0:0:0, 0, notifier);
	$width (posedge BRAMISOCMCLK, 0:0:0, 0, notifier);
	$width (negedge BRAMISOCMCLK, 0:0:0, 0, notifier);
	$width (posedge CPMC405CLOCK, 0:0:0, 0, notifier);
	$width (negedge CPMC405CLOCK, 0:0:0, 0, notifier);
	$width (posedge JTGC405TCK, 0:0:0, 0, notifier);
	$width (negedge JTGC405TCK, 0:0:0, 0, notifier);
	$width (posedge PLBCLK, 0:0:0, 0, notifier);
	$width (negedge PLBCLK, 0:0:0, 0, notifier);
	$period (posedge CPMC405CLOCK, 0:0:0, notifier);

	specparam PATHPULSE$ = 0;

endspecify

endmodule

module FPGA_startup(bus_reset, ghigh_b, gsr, done, gwe, gts_b, shutdown, cclk, por);
   output bus_reset;
   output ghigh_b;
   output gsr;
   output done;
   output gwe;
   output gts_b;
   input  shutdown;
   input  cclk, por;

   reg    bus_reset, abus_reset;
   reg    ghigh_b, aghigh_b;
   reg    gsr, agsr;
   reg    done, adone;
   reg    gwe, agwe;
   reg    gts_b, agts_b;

   reg    [7:0] count;

   always @ (posedge cclk or posedge por) begin
     if(por) count <= {8{1'b0}};
     else if(shutdown && (count > {8{1'b0}})) count = count - 1;
     else if(!shutdown && (count < {8'hFF})) count = count + 1;
   end

   always @ (posedge cclk or posedge por) begin
     if(por) begin
       {bus_reset,ghigh_b,gsr,done,gwe,gts_b} <= 6'b100000;
     end else begin
       {bus_reset,ghigh_b,gsr,done,gwe,gts_b} <= 
                                   {abus_reset,aghigh_b,agsr,adone,agwe,agts_b};
     end
   end

   always @ (count) begin
     // defaults
     
     abus_reset = 1;
     aghigh_b = 0;
     agsr = 0;
     adone = 0;
     agwe = 0;
     agts_b = 0;

     // Trip times are in order for default sequence.
     if(count >= 8'h04) abus_reset = 0;
     if(count == 8'h21 || count == 8'h22) agsr = 1;
     if(count > 8'h26) aghigh_b = 1;
     if(count > 8'h31) adone = 1;
     if(count > 8'h32) agwe = 1;
     if(count > 8'h33) agts_b = 1;
   end
   
endmodule // startup
