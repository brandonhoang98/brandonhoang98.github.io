
/*

FUNCTION	: CONFIG dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module CONFIG ();


endmodule

`endcelldefine
