
/*

FUNCTION	: OPT_OFF dummy simulation module

*/

`timescale  100 ps / 10 ps

`celldefine

module OPT_OFF (I);


    input  I;

endmodule

`endcelldefine
