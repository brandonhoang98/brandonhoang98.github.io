//    Xilinx Proprietary Primitive Cell X_UPAD for Verilog
//
// $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/versclibs/data/X_UPAD.v,v 1.9 2003/01/21 02:38:44 wloo Exp $
//

`timescale 1 ps/1 ps

module X_UPAD (PAD);

  inout PAD;

endmodule
